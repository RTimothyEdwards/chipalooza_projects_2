magic
tech sky130A
magscale 1 2
timestamp 1726321856
<< checkpaint >>
rect 2132 252898 13728 266392
<< metal1 >>
rect 12006 260628 12338 260688
rect 12398 260628 12404 260688
rect 12010 260508 12478 260568
rect 12538 260508 12544 260568
rect 12010 254722 12614 254782
rect 12674 254722 12680 254782
rect 12010 254602 12760 254662
rect 12820 254602 12826 254662
<< via1 >>
rect 12338 260628 12398 260688
rect 12478 260508 12538 260568
rect 12614 254722 12674 254782
rect 12760 254602 12820 254662
<< metal2 >>
rect 4693 259712 5666 261382
rect 12336 260688 12406 260714
rect 12336 260628 12338 260688
rect 12398 260628 12406 260688
rect 12336 252898 12406 260628
rect 12476 260568 12546 260594
rect 12476 260508 12478 260568
rect 12538 260508 12546 260568
rect 12476 252898 12546 260508
rect 12616 254788 12686 254876
rect 12614 254782 12686 254788
rect 12674 254722 12686 254782
rect 12614 254716 12686 254722
rect 12616 252898 12686 254716
rect 12756 254662 12826 254700
rect 12756 254602 12760 254662
rect 12820 254602 12826 254662
rect 12756 252898 12826 254602
<< metal3 >>
rect 8144 266108 13728 266372
rect 11758 260790 13309 261096
rect 11772 259860 13278 260180
rect 11688 253852 13214 254248
rect 2132 253440 5674 253704
rect 8142 253440 13230 253704
use cv3_via2_36cut  cv3_via2_36cut_0
timestamp 1719173892
transform 1 0 -550566 0 1 161218
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_1
timestamp 1719173892
transform 1 0 -547122 0 1 173890
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_2
timestamp 1719173892
transform 1 0 -547114 0 1 161202
box 555256 92202 556228 92502
use switch_array_2  switch_array_2_0
timestamp 1724444975
transform -1 0 11786 0 1 255004
box -328 -1310 7820 11108
<< end >>
