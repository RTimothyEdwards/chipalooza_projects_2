* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_6XHUDR a_n242_n264# a_50_n42# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n242_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6ELFTH a_50_n42# a_n50_n139# w_n308_n339# a_n108_n42#
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n308_n339# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_L7BSKG a_n73_n11# a_n33_n99# a_15_n11# a_n175_n185#
X0 a_15_n11# a_n33_n99# a_n73_n11# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_LGS3BL a_n73_n64# a_n33_n161# a_15_n64# w_n211_n284#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n211_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_64Z3AY a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt rc_osc_level_shifter out_h outb_h in_l dvss inb_l avss dvdd avdd
XXM15 outb_h out_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM16 avdd outb_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM17 avss outb_h avss in_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM18 avss avss out_h inb_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM19 m1_2204_n1198# out_h avdd avdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM7 dvdd in_l inb_l dvdd sky130_fd_pr__pfet_01v8_LGS3BL
XXM8 inb_l dvss in_l dvss sky130_fd_pr__nfet_01v8_64Z3AY
XXM20 m1_2204_n1198# outb_h avdd out_h sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
.ends

.subckt sky130_fd_pr__nfet_01v8_L9WNCD a_15_n19# a_n175_n193# a_n73_n19# a_n33_n107#
X0 a_15_n19# a_n33_n107# a_n73_n19# a_n175_n193# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__3 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__pfet_01v8_856REK a_63_n150# a_15_181# w_n263_n369# a_n81_n247#
+ a_n125_n150#
X0 a_63_n150# a_15_181# a_n33_n150# w_n263_n369# sky130_fd_pr__pfet_01v8 ad=0.465 pd=3.62 as=0.2475 ps=1.83 w=1.5 l=0.15
X1 a_n33_n150# a_n81_n247# a_n125_n150# w_n263_n369# sky130_fd_pr__pfet_01v8 ad=0.2475 pd=1.83 as=0.465 ps=3.62 w=1.5 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF a_2372_n1166# a_3700_n1166# a_n2276_734#
+ a_n1944_n1166# a_n3272_734# a_n3438_n1166# a_n782_n1166# a_1376_n1166# a_1542_734#
+ a_4696_734# a_2704_n1166# a_546_n1166# a_546_734# a_1708_n1166# a_n1114_734# a_n4268_734#
+ a_n118_734# a_2538_734# a_n2110_734# a_n2442_n1166# a_3534_734# a_3202_n1166# a_n1446_n1166#
+ a_4530_734# a_n284_n1166# a_4696_n1166# a_n3106_734# a_2206_n1166# a_n4102_734#
+ a_1874_734# a_n616_n1166# a_n450_734# a_2870_734# a_878_734# a_1210_n1166# a_n1446_734#
+ a_n4766_n1166# a_n2442_734# a_3866_734# a_4198_n1166# a_4862_734# a_878_n1166# a_n118_n1166#
+ a_712_734# a_n3438_734# a_n3770_n1166# a_1708_734# a_n4434_734# a_2704_734# a_4530_n1166#
+ a_n2774_n1166# a_n782_734# a_3700_734# a_n4268_n1166# a_n5062_n1296# a_3534_n1166#
+ a_n1778_n1166# a_n1778_734# a_n2774_734# a_2538_n1166# a_n3770_734# a_n3272_n1166#
+ a_n4600_n1166# a_n948_n1166# a_1044_734# a_380_n1166# a_4198_734# a_4032_n1166#
+ a_n2276_n1166# a_2040_734# a_n3604_n1166# a_n1612_734# a_1542_n1166# a_n4766_734#
+ a_n616_734# a_712_n1166# a_3036_n1166# a_n2608_n1166# a_3036_734# a_n1280_n1166#
+ a_n2608_734# a_4032_734# a_n3604_734# a_n4102_n1166# a_48_734# a_2040_n1166# a_n1612_n1166#
+ a_n4600_734# a_380_734# a_4862_n1166# a_n450_n1166# a_n3106_n1166# a_1044_n1166#
+ a_1376_734# a_214_n1166# a_2372_734# a_3866_n1166# a_n1944_734# a_n948_734# a_n2940_734#
+ a_n2110_n1166# a_3368_734# a_n4932_n1166# a_n1114_n1166# a_1210_734# a_2870_n1166#
+ a_4364_734# a_n3936_734# a_4364_n1166# a_n3936_n1166# a_214_734# a_n4932_734# a_1874_n1166#
+ a_3368_n1166# a_2206_734# a_48_n1166# a_n1280_734# a_n284_734# a_3202_734# a_n2940_n1166#
+ a_n4434_n1166#
X0 a_n4766_734# a_n4766_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X1 a_712_734# a_712_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X2 a_1874_734# a_1874_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X3 a_n3272_734# a_n3272_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X4 a_n1612_734# a_n1612_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X5 a_n3770_734# a_n3770_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X6 a_n782_734# a_n782_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X7 a_n2276_734# a_n2276_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X8 a_n118_734# a_n118_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X9 a_4696_734# a_4696_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X10 a_n4434_734# a_n4434_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X11 a_1542_734# a_1542_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X12 a_n1280_734# a_n1280_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X13 a_3700_734# a_3700_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X14 a_n3438_734# a_n3438_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X15 a_4364_734# a_4364_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X16 a_n948_734# a_n948_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X17 a_2704_734# a_2704_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X18 a_n4102_734# a_n4102_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X19 a_1210_734# a_1210_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X20 a_1708_734# a_1708_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X21 a_3368_734# a_3368_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X22 a_n3106_734# a_n3106_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X23 a_n2774_734# a_n2774_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X24 a_n616_734# a_n616_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X25 a_380_734# a_380_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X26 a_4032_734# a_4032_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X27 a_n2110_734# a_n2110_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X28 a_n4932_734# a_n4932_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X29 a_878_734# a_878_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X30 a_3036_734# a_3036_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X31 a_n1778_734# a_n1778_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X32 a_n3936_734# a_n3936_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X33 a_n2442_734# a_n2442_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X34 a_4862_734# a_4862_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X35 a_n4600_734# a_n4600_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X36 a_n2940_734# a_n2940_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X37 a_546_734# a_546_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X38 a_n1446_734# a_n1446_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X39 a_3866_734# a_3866_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X40 a_n3604_734# a_n3604_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X41 a_2372_734# a_2372_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X42 a_4530_734# a_4530_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X43 a_n4268_734# a_n4268_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X44 a_214_734# a_214_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X45 a_1376_734# a_1376_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X46 a_n2608_734# a_n2608_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X47 a_n1114_734# a_n1114_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X48 a_2040_734# a_2040_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X49 a_3534_734# a_3534_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X50 a_n284_734# a_n284_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X51 a_2538_734# a_2538_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X52 a_4198_734# a_4198_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X53 a_1044_734# a_1044_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X54 a_3202_734# a_3202_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X55 a_n1944_734# a_n1944_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X56 a_n450_734# a_n450_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X57 a_48_734# a_48_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X58 a_2206_734# a_2206_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
X59 a_2870_734# a_2870_n1166# a_n5062_n1296# sky130_fd_pr__res_xhigh_po_0p35 l=7.5
.ends

.subckt sky130_fd_pr__pfet_01v8_2Z69BZ w_n211_n226# a_n73_n6# a_15_n6# a_n33_n103#
X0 a_15_n6# a_n33_n103# a_n73_n6# w_n211_n226# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_T537S5 a_n50_n223# w_n308_n423# a_50_n126# a_n108_n126#
X0 a_50_n126# a_n50_n223# a_n108_n126# w_n308_n423# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.5
.ends

.subckt sky130_ef_ip__rc_osc_16M avdd dvdd ena dout dvss avss
XXM12 avss m1_6428_4585# avss m1_2993_5163# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM34 avdd m1_1507_5567# avdd m1_1507_5567# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM23 avss m1_5241_4130# m1_513_6590# rc_osc_level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM35 dout rc_osc_level_shifter_0/inb_l dvss dvss sky130_fd_pr__nfet_01v8_L7BSKG
XXM13 avss m1_6642_4785# m1_6428_4585# ena sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM25 avdd m1_1507_5567# avdd m1_3601_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM24 avdd m1_1507_5567# avdd m1_2985_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM36 avss m1_2561_4188# m1_1507_5567# rc_osc_level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM26 avdd m1_1507_5567# avdd m1_4217_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM15 m1_2993_5163# m1_4789_4781# avdd m1_5449_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM16 avss m1_2993_5163# m1_5128_4639# m1_4789_4781# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM27 avss m1_4016_4639# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM17 avdd m1_1507_5567# avdd m1_4833_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM28 avss m1_3460_4639# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xrc_osc_level_shifter_0 rc_osc_level_shifter_0/out_h rc_osc_level_shifter_0/outb_h
+ ena dvss rc_osc_level_shifter_0/inb_l avss dvdd avdd rc_osc_level_shifter
XXM18 avdd m1_1507_5567# avdd m1_1507_5567# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM29 avss m1_2904_4639# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM19 avss m1_5128_4639# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM1 avss m1_3128_4787# m1_2904_4639# m1_2993_5163# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM2 m1_3128_4787# m1_2993_5163# avdd m1_2985_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM3 m1_3679_4781# m1_3128_4787# avdd m1_3601_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM4 avss m1_3679_4781# m1_3460_4639# m1_3128_4787# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xsky130_fd_pr__nfet_01v8_L9WNCD_0 dout dvss dvss m1_6642_4785# sky130_fd_pr__nfet_01v8_L9WNCD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__3
XXM7 m1_4789_4781# m1_4235_4789# avdd m1_4833_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM9 m1_4235_4789# m1_3679_4781# avdd m1_4217_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM8 avss m1_4789_4781# m1_4572_4639# m1_4235_4789# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_0 avdd m1_1507_5567# avdd m1_1507_5567# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__pfet_01v8_856REK_0 dout rc_osc_level_shifter_0/inb_l dvdd m1_6642_4785#
+ dvdd sky130_fd_pr__pfet_01v8_856REK
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_1 avdd m1_1507_5567# avdd m1_1507_5567# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_0 m1_7838_1218# m1_9166_1218# m1_3024_3118#
+ m1_3522_1218# m1_2028_3118# m1_1862_1218# m1_4518_1218# m1_6842_1218# m1_7008_3118#
+ m1_9996_3118# m1_8170_1218# m1_5846_1218# m1_6012_3118# m1_7174_1218# m1_4352_3118#
+ m1_1032_3118# m1_5348_3118# m1_8004_3118# m1_3356_3118# m1_2858_1218# m1_9000_3118#
+ m1_8502_1218# m1_3854_1218# m1_9996_3118# m1_5182_1218# m1_10162_1218# m1_2360_3118#
+ m1_7506_1218# m1_1364_3118# m1_7340_3118# m1_4850_1218# m1_5016_3118# m1_8336_3118#
+ m1_6344_3118# m1_6510_1218# m1_4020_3118# m1_534_1218# m1_3024_3118# m1_9332_3118#
+ m1_9498_1218# m1_9378_4056# m1_6178_1218# m1_5182_1218# m1_6012_3118# m1_2028_3118#
+ m1_1530_1218# m1_7008_3118# m1_1032_3118# m1_8004_3118# m1_9830_1218# m1_2526_1218#
+ m1_4684_3118# m1_9000_3118# m1_1198_1218# avss m1_8834_1218# m1_3522_1218# m1_3688_3118#
+ m1_2692_3118# m1_7838_1218# m1_1696_3118# m1_2194_1218# m1_866_1218# m1_4518_1218#
+ m1_6344_3118# m1_5846_1218# m1_9664_3118# m1_9498_1218# m1_3190_1218# m1_7340_3118#
+ m1_1862_1218# m1_3688_3118# m1_6842_1218# m1_700_3118# m1_4684_3118# m1_6178_1218#
+ m1_8502_1218# m1_2858_1218# m1_8336_3118# m1_4186_1218# m1_2692_3118# m1_9332_3118#
+ m1_1696_3118# m1_1198_1218# m1_5348_3118# m1_7506_1218# m1_3854_1218# m1_700_3118#
+ m1_5680_3118# m1_10162_1218# m1_4850_1218# m1_2194_1218# m1_6510_1218# m1_6676_3118#
+ m1_5514_1218# m1_7672_3118# m1_9166_1218# m1_3356_3118# m1_4352_3118# m1_2360_3118#
+ m1_3190_1218# m1_8668_3118# m1_534_1218# m1_4186_1218# m1_6676_3118# m1_8170_1218#
+ m1_9664_3118# m1_1364_3118# m1_9830_1218# m1_1530_1218# m1_5680_3118# avdd m1_7174_1218#
+ m1_8834_1218# m1_7672_3118# m1_5514_1218# m1_4020_3118# m1_5016_3118# m1_8668_3118#
+ m1_2526_1218# m1_866_1218# sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF
Xsky130_fd_pr__res_xhigh_po_0p35_NVJ5PF_1 m1_7652_7168# m1_8980_7168# m1_3170_9068#
+ m1_3336_7168# m1_2174_9068# m1_2008_7168# m1_4664_7168# m1_6656_7168# m1_6822_9068#
+ m1_10142_9068# m1_7984_7168# m1_5992_7168# m1_5826_9068# m1_6988_7168# m1_4166_9068#
+ m1_1178_9068# m1_5162_9068# m1_7818_9068# m1_3170_9068# m1_3004_7168# m1_8814_9068#
+ m1_8648_7168# m1_4000_7168# m1_9810_9068# m1_4996_7168# m1_9976_7168# m1_2174_9068#
+ m1_7652_7168# m1_1178_9068# m1_7154_9068# m1_4664_7168# m1_4830_9068# m1_8150_9068#
+ m1_6158_9068# m1_6656_7168# m1_3834_9068# m1_680_7168# avdd m1_9146_9068# m1_9644_7168#
+ m1_10142_9068# m1_6324_7168# m1_5328_7168# m1_6158_9068# m1_1842_9068# m1_1676_7168#
+ m1_7154_9068# m1_846_9068# m1_8150_9068# m1_9976_7168# m1_2672_7168# m1_4498_9068#
+ m1_9146_9068# m1_1012_7168# avss m1_8980_7168# m1_3668_7168# m1_3502_9068# m1_2506_9068#
+ m1_7984_7168# m1_1510_9068# m1_2008_7168# m1_680_7168# m1_4332_7168# m1_6490_9068#
+ m1_5660_7168# m1_9478_9068# m1_9312_7168# m1_3004_7168# m1_7486_9068# m1_1676_7168#
+ m1_3834_9068# m1_6988_7168# m1_514_9068# m1_4830_9068# m1_5992_7168# m1_8316_7168#
+ m1_2672_7168# m1_8482_9068# m1_4000_7168# avdd m1_9478_9068# m1_1842_9068# m1_1344_7168#
+ m1_5494_9068# m1_7320_7168# m1_3668_7168# m1_846_9068# m1_5826_9068# m1_9378_4056#
+ m1_4996_7168# m1_2340_7168# m1_6324_7168# m1_6822_9068# m1_5660_7168# m1_7818_9068#
+ m1_9312_7168# m1_3502_9068# m1_4498_9068# m1_2506_9068# m1_3336_7168# m1_8814_9068#
+ m1_513_6590# m1_4332_7168# m1_6490_9068# m1_8316_7168# m1_9810_9068# m1_1510_9068#
+ m1_9644_7168# m1_1344_7168# m1_5494_9068# m1_514_9068# m1_7320_7168# m1_8648_7168#
+ m1_7486_9068# m1_5328_7168# m1_4166_9068# m1_5162_9068# m1_8482_9068# m1_2340_7168#
+ m1_1012_7168# sky130_fd_pr__res_xhigh_po_0p35_NVJ5PF
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_2 m1_1507_5567# m1_1507_5567# avdd avdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_3 avdd rc_osc_level_shifter_0/out_h avdd m1_1507_5567#
+ sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__pfet_01v8_2Z69BZ_0 dvdd m1_6642_4785# dvdd ena sky130_fd_pr__pfet_01v8_2Z69BZ
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_5 avdd m1_1507_5567# avdd m1_5449_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__pfet_g5v0d10v5_6ELFTH_4 m1_1507_5567# m1_1507_5567# avdd avdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xsky130_fd_pr__pfet_g5v0d10v5_T537S5_0 m1_2993_5163# avdd m1_6642_4785# dvdd sky130_fd_pr__pfet_g5v0d10v5_T537S5
XXM30 avss m1_2561_4188# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM20 avss m1_4572_4639# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM10 avss m1_4235_4789# m1_4016_4639# m1_3679_4781# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM21 avss m1_5241_4130# avss m1_5241_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM33 avss m1_5241_4130# avss rc_osc_level_shifter_0/outb_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WQT6C6 a_1235_n700# a_3447_n700# a_5659_n700#
+ a_n287_n788# a_761_n700# a_n4079_n788# a_819_n788# a_2657_n700# a_4869_n700# a_5185_n700#
+ a_n1077_n788# a_n3289_n788# a_1867_n700# a_2183_n700# a_345_n788# a_4395_n700# a_n29_n700#
+ a_n2499_n788# a_1393_n700# a_n919_n788# a_6607_n700# a_977_n788# a_n5027_n788# a_3605_n700#
+ a_5817_n700# a_n445_n788# a_3189_n788# a_n187_n700# a_6133_n700# a_n1709_n788# a_n2025_n788#
+ a_n4237_n788# a_2815_n700# a_n6449_n788# a_3131_n700# a_5343_n700# a_2399_n788#
+ a_n1235_n788# a_n3447_n788# a_n5659_n788# a_n3189_n700# a_2341_n700# a_4553_n700#
+ a_503_n788# a_6765_n700# a_n2657_n788# a_n4869_n788# a_n5185_n788# a_n2399_n700#
+ a_1551_n700# a_3763_n700# a_5975_n700# a_1609_n788# a_6291_n700# a_n1867_n788# a_6349_n788#
+ a_n819_n700# a_4137_n788# a_n2183_n788# a_n4395_n788# a_2973_n700# a_n603_n788#
+ a_3347_n788# a_1135_n788# a_n7124_n700# a_n345_n700# a_5559_n788# a_n1393_n788#
+ a_n1609_n700# a_n6607_n788# a_661_n788# a_n6349_n700# a_n4137_n700# a_5501_n700#
+ a_4769_n788# a_2557_n788# a_5085_n788# a_n3605_n788# a_n5817_n788# a_n3347_n700#
+ a_n1135_n700# a_n6133_n788# a_n5559_n700# a_4711_n700# a_6923_n700# a_3979_n788#
+ a_1767_n788# a_n977_n700# a_4295_n788# a_2083_n788# a_n2815_n788# a_n3131_n788#
+ a_n5343_n788# a_n4769_n700# a_n2557_n700# a_3921_n700# a_n5085_n700# a_1293_n788#
+ a_n761_n788# a_6507_n788# a_n2341_n788# a_n3979_n700# a_n1767_n700# a_n4553_n788#
+ a_n6765_n788# a_n4295_n700# a_n2083_n700# a_5717_n788# a_3505_n788# a_6033_n788#
+ a_n503_n700# a_n1551_n788# a_n3763_n788# a_n5975_n788# a_n1293_n700# a_129_n700#
+ a_n6291_n788# a_n6507_n700# a_2715_n788# a_4927_n788# a_3031_n788# a_n2973_n788#
+ a_5243_n788# a_n5717_n700# a_n3505_n700# a_n6033_n700# a_1925_n788# a_4453_n788#
+ a_2241_n788# a_6665_n788# a_n2715_n700# a_n5501_n788# a_n4927_n700# a_n3031_n700#
+ a_n5243_n700# a_1451_n788# a_5875_n788# a_n661_n700# a_3663_n788# a_6191_n788# a_287_n700#
+ a_n4711_n788# a_n1925_n700# a_n6923_n788# a_n4453_n700# a_n2241_n700# a_n6665_n700#
+ a_2873_n788# a_n3921_n788# a_n1451_n700# a_n5875_n700# a_n3663_n700# a_n6191_n700#
+ a_5401_n788# a_n2873_n700# a_6823_n788# a_4611_n788# a_919_n700# a_n5401_n700# a_3821_n788#
+ a_445_n700# a_n6823_n700# a_n4611_n700# a_n3821_n700# a_4079_n700# a_1077_n700#
+ a_3289_n700# a_29_n788# a_2499_n700# a_n6981_n700# a_n129_n788# a_603_n700# a_187_n788#
+ a_5027_n700# a_1709_n700# a_2025_n700# a_4237_n700# a_6449_n700#
X0 a_n6349_n700# a_n6449_n788# a_n6507_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X1 a_n5875_n700# a_n5975_n788# a_n6033_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X2 a_n3505_n700# a_n3605_n788# a_n3663_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X3 a_3605_n700# a_3505_n788# a_3447_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X4 a_5975_n700# a_5875_n788# a_5817_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X5 a_6449_n700# a_6349_n788# a_6291_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X6 a_n6191_n700# a_n6291_n788# a_n6349_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X7 a_n977_n700# a_n1077_n788# a_n1135_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X8 a_6291_n700# a_6191_n788# a_6133_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X9 a_n503_n700# a_n603_n788# a_n661_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X10 a_1077_n700# a_977_n788# a_919_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X11 a_n5401_n700# a_n5501_n788# a_n5559_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X12 a_n2557_n700# a_n2657_n788# a_n2715_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X13 a_2657_n700# a_2557_n788# a_2499_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X14 a_5501_n700# a_5401_n788# a_5343_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X15 a_n4927_n700# a_n5027_n788# a_n5085_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X16 a_n4453_n700# a_n4553_n788# a_n4611_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X17 a_n29_n700# a_n129_n788# a_n187_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X18 a_603_n700# a_503_n788# a_445_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X19 a_4553_n700# a_4453_n788# a_4395_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X20 a_n6507_n700# a_n6607_n788# a_n6665_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X21 a_6607_n700# a_6507_n788# a_6449_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X22 a_n3979_n700# a_n4079_n788# a_n4137_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X23 a_n1135_n700# a_n1235_n788# a_n1293_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X24 a_1235_n700# a_1135_n788# a_1077_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X25 a_5659_n700# a_5559_n788# a_5501_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X26 a_n5559_n700# a_n5659_n788# a_n5717_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X27 a_n2715_n700# a_n2815_n788# a_n2873_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X28 a_2815_n700# a_2715_n788# a_2657_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X29 a_n3031_n700# a_n3131_n788# a_n3189_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X30 a_3131_n700# a_3031_n788# a_2973_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X31 a_n4611_n700# a_n4711_n788# a_n4769_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X32 a_n1767_n700# a_n1867_n788# a_n1925_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X33 a_1867_n700# a_1767_n788# a_1709_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X34 a_4711_n700# a_4611_n788# a_4553_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X35 a_2183_n700# a_2083_n788# a_2025_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X36 a_n2083_n700# a_n2183_n788# a_n2241_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X37 a_n4137_n700# a_n4237_n788# a_n4295_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X38 a_n3663_n700# a_n3763_n788# a_n3821_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X39 a_3763_n700# a_3663_n788# a_3605_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X40 a_4237_n700# a_4137_n788# a_4079_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X41 a_n819_n700# a_n919_n788# a_n977_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X42 a_n5717_n700# a_n5817_n788# a_n5875_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X43 a_n661_n700# a_n761_n788# a_n819_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X44 a_5817_n700# a_5717_n788# a_5659_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X45 a_n6033_n700# a_n6133_n788# a_n6191_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X46 a_n3189_n700# a_n3289_n788# a_n3347_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X47 a_3289_n700# a_3189_n788# a_3131_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X48 a_6133_n700# a_6033_n788# a_5975_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X49 a_n4769_n700# a_n4869_n788# a_n4927_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X50 a_919_n700# a_819_n788# a_761_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X51 a_2025_n700# a_1925_n788# a_1867_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X52 a_4869_n700# a_4769_n788# a_4711_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X53 a_n5085_n700# a_n5185_n788# a_n5243_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X54 a_n187_n700# a_n287_n788# a_n345_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X55 a_761_n700# a_661_n788# a_603_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X56 a_5185_n700# a_5085_n788# a_5027_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X57 a_n2241_n700# a_n2341_n788# a_n2399_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X58 a_2341_n700# a_2241_n788# a_2183_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X59 a_n6665_n700# a_n6765_n788# a_n6823_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X60 a_n3821_n700# a_n3921_n788# a_n3979_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X61 a_287_n700# a_187_n788# a_129_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X62 a_3921_n700# a_3821_n788# a_3763_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X63 a_6765_n700# a_6665_n788# a_6607_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X64 a_n1293_n700# a_n1393_n788# a_n1451_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X65 a_1393_n700# a_1293_n788# a_1235_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X66 a_n3347_n700# a_n3447_n788# a_n3505_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X67 a_n2873_n700# a_n2973_n788# a_n3031_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X68 a_2973_n700# a_2873_n788# a_2815_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X69 a_3447_n700# a_3347_n788# a_3289_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X70 a_5027_n700# a_4927_n788# a_4869_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X71 a_n345_n700# a_n445_n788# a_n503_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X72 a_2499_n700# a_2399_n788# a_2341_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X73 a_5343_n700# a_5243_n788# a_5185_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X74 a_n5243_n700# a_n5343_n788# a_n5401_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X75 a_n2399_n700# a_n2499_n788# a_n2557_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X76 a_n6823_n700# a_n6923_n788# a_n6981_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X77 a_n1609_n700# a_n1709_n788# a_n1767_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X78 a_129_n700# a_29_n788# a_n29_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X79 a_1709_n700# a_1609_n788# a_1551_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X80 a_4079_n700# a_3979_n788# a_3921_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X81 a_6923_n700# a_6823_n788# a_6765_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X82 a_n4295_n700# a_n4395_n788# a_n4453_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X83 a_n1925_n700# a_n2025_n788# a_n2083_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X84 a_n1451_n700# a_n1551_n788# a_n1609_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X85 a_445_n700# a_345_n788# a_287_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X86 a_1551_n700# a_1451_n788# a_1393_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X87 a_4395_n700# a_4295_n788# a_4237_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7WGKBW a_5875_n1597# a_5343_n1500# a_n761_n1597#
+ a_3131_n1500# a_5817_n1500# a_3663_n1597# a_187_n1597# a_129_n1500# a_3605_n1500#
+ a_1451_n1597# a_1925_n1597# a_n2399_n1500# a_n6133_n1597# a_5185_n1500# a_661_n1597#
+ a_n6607_n1597# a_5659_n1500# a_603_n1500# a_3447_n1500# a_3979_n1597# a_1293_n1597#
+ a_n2873_n1500# a_1767_n1597# a_1235_n1500# a_1709_n1500# a_n6449_n1597# a_3921_n1500#
+ a_977_n1597# a_445_n1500# a_n4237_n1597# a_919_n1500# a_3289_n1500# a_n2025_n1597#
+ a_6033_n1597# a_1077_n1500# a_6507_n1597# a_n6923_n1597# a_5975_n1500# a_n5401_n1500#
+ a_n4711_n1597# a_287_n1500# a_3763_n1500# a_n4079_n1597# a_1551_n1500# a_n6291_n1597#
+ a_6349_n1597# a_n6765_n1597# a_761_n1500# a_n5243_n1500# a_n29_n1500# a_4137_n1597#
+ a_n4553_n1597# a_n5717_n1500# a_n3031_n1500# a_n2341_n1597# a_1393_n1500# a_n3505_n1500#
+ a_n2815_n1597# a_6823_n1597# a_1867_n1500# a_4611_n1597# a_n5085_n1500# a_n4395_n1597#
+ a_n5559_n1500# a_6191_n1597# a_n2183_n1597# a_n4869_n1597# a_n3347_n1500# a_6665_n1597#
+ a_6133_n1500# a_n2657_n1597# a_n1135_n1500# a_6607_n1500# a_4453_n1597# a_n1609_n1500#
+ a_4927_n1597# a_n503_n1500# a_2241_n1597# a_n3821_n1500# a_2715_n1597# a_n3189_n1500#
+ a_n2499_n1597# a_6449_n1500# a_4295_n1597# a_n5875_n1500# a_4237_n1500# a_4769_n1597#
+ a_2083_n1597# a_n345_n1500# a_n3663_n1500# a_2025_n1500# a_2557_n1597# a_n2973_n1597#
+ a_n819_n1500# a_n1451_n1500# a_6923_n1500# a_n1925_n1500# a_4711_n1500# a_29_n1597#
+ a_n5027_n1597# a_4079_n1500# a_n187_n1500# a_2399_n1597# a_6291_n1500# a_n3979_n1500#
+ a_n1293_n1500# a_6765_n1500# a_n1767_n1500# a_n5501_n1597# a_4553_n1500# a_n661_n1500#
+ a_2341_n1500# a_2873_n1597# a_2815_n1500# a_n6033_n1500# a_n5343_n1597# a_n6507_n1500#
+ a_4395_n1500# a_n3131_n1597# a_n5817_n1597# a_n977_n1500# a_2183_n1500# a_4869_n1500#
+ a_n3605_n1597# a_2657_n1500# a_5401_n1597# a_n5185_n1597# a_n6349_n1500# a_n5659_n1597#
+ a_n129_n1597# a_n4137_n1500# a_n3447_n1597# a_2499_n1500# a_5243_n1597# a_n1235_n1597#
+ a_n1709_n1597# a_n6823_n1500# a_5717_n1597# a_3031_n1597# a_n603_n1597# a_n4611_n1500#
+ a_3505_n1597# a_n3921_n1597# a_2973_n1500# a_n3289_n1597# a_n1077_n1597# a_n6191_n1500#
+ a_5085_n1597# w_n7017_n1600# a_n6665_n1500# a_5027_n1500# a_5559_n1597# a_503_n1597#
+ a_n5975_n1597# a_n445_n1597# a_n4453_n1500# a_3347_n1597# a_n3763_n1597# a_n919_n1597#
+ a_n4927_n1500# a_n2241_n1500# a_1135_n1597# a_n1551_n1597# a_n2715_n1500# a_1609_n1597#
+ a_5501_n1500# a_3821_n1597# a_345_n1597# a_n287_n1597# a_n4295_n1500# a_3189_n1597#
+ a_819_n1597# a_n4769_n1500# a_n2083_n1500# a_n1393_n1597# a_n6981_n1500# a_n2557_n1500#
+ a_n1867_n1597#
X0 a_n6033_n1500# a_n6133_n1597# a_n6191_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X1 a_n819_n1500# a_n919_n1597# a_n977_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X2 a_n6191_n1500# a_n6291_n1597# a_n6349_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X3 a_n977_n1500# a_n1077_n1597# a_n1135_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X4 a_2973_n1500# a_2873_n1597# a_2815_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X5 a_n6507_n1500# a_n6607_n1597# a_n6665_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X6 a_1235_n1500# a_1135_n1597# a_1077_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X7 a_1393_n1500# a_1293_n1597# a_1235_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X8 a_4079_n1500# a_3979_n1597# a_3921_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X9 a_n6665_n1500# a_n6765_n1597# a_n6823_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X10 a_603_n1500# a_503_n1597# a_445_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X11 a_1709_n1500# a_1609_n1597# a_1551_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X12 a_n4927_n1500# a_n5027_n1597# a_n5085_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X13 a_761_n1500# a_661_n1597# a_603_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X14 a_6923_n1500# a_6823_n1597# a_6765_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=0.5
X15 a_n5085_n1500# a_n5185_n1597# a_n5243_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X16 a_n4453_n1500# a_n4553_n1597# a_n4611_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X17 a_n3821_n1500# a_n3921_n1597# a_n3979_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X18 a_1867_n1500# a_1767_n1597# a_1709_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X19 a_2499_n1500# a_2399_n1597# a_2341_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X20 a_4711_n1500# a_4611_n1597# a_4553_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X21 a_5343_n1500# a_5243_n1597# a_5185_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X22 a_n2241_n1500# a_n2341_n1597# a_n2399_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X23 a_n5559_n1500# a_n5659_n1597# a_n5717_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X24 a_3131_n1500# a_3031_n1597# a_2973_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X25 a_n503_n1500# a_n603_n1597# a_n661_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X26 a_5817_n1500# a_5717_n1597# a_5659_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X27 a_6449_n1500# a_6349_n1597# a_6291_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X28 a_n3347_n1500# a_n3447_n1597# a_n3505_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X29 a_n2715_n1500# a_n2815_n1597# a_n2873_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X30 a_287_n1500# a_187_n1597# a_129_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X31 a_5975_n1500# a_5875_n1597# a_5817_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X32 a_n3979_n1500# a_n4079_n1597# a_n4137_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X33 a_n2873_n1500# a_n2973_n1597# a_n3031_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X34 a_n661_n1500# a_n761_n1597# a_n819_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X35 a_3605_n1500# a_3505_n1597# a_3447_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X36 a_4237_n1500# a_4137_n1597# a_4079_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X37 a_n1135_n1500# a_n1235_n1597# a_n1293_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X38 a_3763_n1500# a_3663_n1597# a_3605_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X39 a_4395_n1500# a_4295_n1597# a_4237_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X40 a_n1293_n1500# a_n1393_n1597# a_n1451_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X41 a_n6823_n1500# a_n6923_n1597# a_n6981_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=0.5
X42 a_n1609_n1500# a_n1709_n1597# a_n1767_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X43 a_n29_n1500# a_n129_n1597# a_n187_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X44 a_1551_n1500# a_1451_n1597# a_1393_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X45 a_2183_n1500# a_2083_n1597# a_2025_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X46 a_4869_n1500# a_4769_n1597# a_4711_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X47 a_n1767_n1500# a_n1867_n1597# a_n1925_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X48 a_n187_n1500# a_n287_n1597# a_n345_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X49 a_n4611_n1500# a_n4711_n1597# a_n4769_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X50 a_n2399_n1500# a_n2499_n1597# a_n2557_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X51 a_2025_n1500# a_1925_n1597# a_1867_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X52 a_n5243_n1500# a_n5343_n1597# a_n5401_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X53 a_2657_n1500# a_2557_n1597# a_2499_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X54 a_3289_n1500# a_3189_n1597# a_3131_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X55 a_5501_n1500# a_5401_n1597# a_5343_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X56 a_6133_n1500# a_6033_n1597# a_5975_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X57 a_n5717_n1500# a_n5817_n1597# a_n5875_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X58 a_n3031_n1500# a_n3131_n1597# a_n3189_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X59 a_129_n1500# a_29_n1597# a_n29_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X60 a_n6349_n1500# a_n6449_n1597# a_n6507_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X61 a_6291_n1500# a_6191_n1597# a_6133_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X62 a_n5875_n1500# a_n5975_n1597# a_n6033_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X63 a_445_n1500# a_345_n1597# a_287_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X64 a_6607_n1500# a_6507_n1597# a_6449_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X65 a_n4137_n1500# a_n4237_n1597# a_n4295_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X66 a_n3505_n1500# a_n3605_n1597# a_n3663_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X67 a_6765_n1500# a_6665_n1597# a_6607_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X68 a_n3663_n1500# a_n3763_n1597# a_n3821_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X69 a_n4295_n1500# a_n4395_n1597# a_n4453_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X70 a_n1925_n1500# a_n2025_n1597# a_n2083_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X71 a_919_n1500# a_819_n1597# a_761_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X72 a_3921_n1500# a_3821_n1597# a_3763_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X73 a_4553_n1500# a_4453_n1597# a_4395_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X74 a_n1451_n1500# a_n1551_n1597# a_n1609_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X75 a_1077_n1500# a_977_n1597# a_919_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X76 a_5185_n1500# a_5085_n1597# a_5027_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X77 a_n4769_n1500# a_n4869_n1597# a_n4927_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X78 a_n2083_n1500# a_n2183_n1597# a_n2241_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X79 a_2341_n1500# a_2241_n1597# a_2183_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X80 a_5027_n1500# a_4927_n1597# a_4869_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X81 a_5659_n1500# a_5559_n1597# a_5501_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X82 a_n2557_n1500# a_n2657_n1597# a_n2715_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X83 a_n345_n1500# a_n445_n1597# a_n503_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X84 a_n5401_n1500# a_n5501_n1597# a_n5559_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X85 a_n3189_n1500# a_n3289_n1597# a_n3347_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X86 a_2815_n1500# a_2715_n1597# a_2657_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X87 a_3447_n1500# a_3347_n1597# a_3289_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3BH9ZH a_n345_n200# a_129_n200# a_287_n200# a_428_n196#
+ a_29_n288# a_n129_n288# a_187_n288# a_n287_n288# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n288# a_n29_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n288# a_n187_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RTDP6L a_n29_n400# w_n381_n500# a_n187_n400#
+ a_n345_n400# a_29_n497# a_n129_n497# a_187_n497# a_129_n400# a_n287_n497# a_287_n400#
X0 a_n29_n400# a_n129_n497# a_n187_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n187_n400# a_n287_n497# a_n345_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2 a_287_n400# a_187_n497# a_129_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_129_n400# a_29_n497# a_n29_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt gate_drive in_m in_p out vdd vss vsub
Xxm1 vss vss vss li_n2466_n1927# out li_n5626_n1927# li_n2466_n1927# out out out li_n2466_n1927#
+ li_n5626_n1927# vss vss li_n2466_n1927# vss vss li_n2466_n1927# out li_n2466_n1927#
+ vss li_n2466_n1927# li_n5626_n1927# out out li_n2466_n1927# li_n2466_n1927# out
+ out li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# vss li_n6574_n1927# vss vss
+ li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# li_n5626_n1927# vss out out li_n2466_n1927#
+ out li_n5626_n1927# li_n5626_n1927# li_n5626_n1927# out vss vss vss li_n2466_n1927#
+ vss li_n2466_n1927# li_n2466_n1927# out li_n2466_n1927# li_n2466_n1927# li_n5626_n1927#
+ out li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# vss vss li_n2466_n1927# li_n2466_n1927#
+ vss li_n6574_n1927# li_n2466_n1927# vss vss out li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n5626_n1927# li_n6574_n1927# li_n2466_n1927# out li_n6574_n1927#
+ li_n2466_n1927# vss vss li_n2466_n1927# li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n5626_n1927# li_n5626_n1927# vss vss out vss li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# out li_n5626_n1927#
+ li_n7839_364# li_n2466_n1927# out li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# li_n6574_n1927# vss out li_n6574_n1927# li_n5626_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# li_n2466_n1927#
+ vss vss vss li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927# vss li_n5626_n1927# vss li_n7839_364#
+ vss vss vss li_n2466_n1927# li_n5626_n1927# out li_n5626_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927# vss vss li_n2466_n1927#
+ out li_n6574_n1927# li_n2466_n1927# vss vss out out li_n2466_n1927# vss vss li_n2466_n1927#
+ vss li_n2466_n1927# vss out out out out sky130_fd_pr__nfet_g5v0d10v5_WQT6C6
Xxm2 li_n2466_n1927# vdd li_n2466_n1927# vdd out li_n2466_n1927# li_n2466_n1927# out
+ out li_n2466_n1927# li_n2466_n1927# out li_n6574_n1927# out li_n2466_n1927# li_n6574_n1927#
+ vdd vdd vdd li_n2466_n1927# li_n2466_n1927# vdd li_n2466_n1927# vdd out li_n6574_n1927#
+ out li_n2466_n1927# out li_n5626_n1927# vdd out li_n2466_n1927# li_n2466_n1927#
+ out li_n2466_n1927# li_n7839_364# vdd vdd li_n5626_n1927# vdd vdd li_n5626_n1927#
+ vdd li_n6574_n1927# li_n2466_n1927# li_n7839_364# out li_n2466_n1927# vdd li_n2466_n1927#
+ li_n5626_n1927# vdd li_n2466_n1927# li_n2466_n1927# out vdd li_n5626_n1927# li_n2466_n1927#
+ vdd li_n2466_n1927# vdd li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# out li_n5626_n1927# out vdd li_n2466_n1927#
+ vdd li_n2466_n1927# out li_n2466_n1927# vdd li_n2466_n1927# vdd li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# out li_n2466_n1927# li_n2466_n1927# vdd li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# out out vdd vdd vdd li_n2466_n1927# li_n5626_n1927#
+ vdd out li_n2466_n1927# vdd li_n2466_n1927# vdd out out li_n5626_n1927# out vdd
+ out li_n2466_n1927# vdd vdd li_n5626_n1927# li_n5626_n1927# vdd li_n5626_n1927#
+ li_n6574_n1927# vdd vdd out li_n5626_n1927# out li_n2466_n1927# li_n5626_n1927#
+ vdd li_n5626_n1927# li_n2466_n1927# vdd li_n5626_n1927# vdd li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n6574_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# out li_n5626_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# vdd vdd vdd li_n2466_n1927# li_n2466_n1927# li_n6574_n1927#
+ li_n2466_n1927# vdd li_n2466_n1927# li_n5626_n1927# li_n2466_n1927# li_n2466_n1927#
+ vdd li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# out li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ vdd out li_n2466_n1927# vdd vdd li_n2466_n1927# sky130_fd_pr__pfet_g5v0d10v5_7WGKBW
Xxm3 vss li_n7839_364# vss vss in_m in_p in_m in_p vss li_n7529_279# sky130_fd_pr__nfet_g5v0d10v5_3BH9ZH
Xxm4 vdd vdd li_n7529_279# vdd li_n7529_279# li_n7839_364# li_n7529_279# li_n7839_364#
+ li_n7839_364# vdd sky130_fd_pr__pfet_g5v0d10v5_RTDP6L
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt pmos_waffle_48x48 dw_n11050_n11060# w_n10844_n10854# a_n50_n50# a_112_3350#
+ a_112_1150#
X0 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X16 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X18 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X19 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X20 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X21 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X22 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X23 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X25 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X26 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X27 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X28 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X30 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X31 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X32 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X33 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X34 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X35 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X36 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X37 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X38 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X39 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X40 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X42 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X43 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X44 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X45 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X46 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X47 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X48 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X49 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X50 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X51 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X52 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X53 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X54 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X55 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X56 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X57 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X58 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X60 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X61 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X62 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X63 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X64 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X65 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X66 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X67 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X68 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X69 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X70 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X71 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X72 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X74 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X75 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X76 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X77 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X78 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X79 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X80 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X81 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X82 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X83 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X84 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X85 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X86 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X87 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X88 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X89 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X90 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X91 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X92 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X93 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X94 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X95 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X96 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X97 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X98 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X99 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X100 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X101 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X104 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X105 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X113 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X115 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X116 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X118 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X119 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X120 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X123 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X136 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X141 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X148 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X149 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X151 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X152 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X157 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X160 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X167 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X168 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X171 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X173 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X182 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X186 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X187 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X188 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X192 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X193 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X196 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X207 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X213 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X214 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X216 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X218 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X224 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X230 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X232 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X233 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X235 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X236 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X238 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X247 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X253 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X255 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X257 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X261 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X263 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X266 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X268 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X270 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X276 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X278 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X279 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X285 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X288 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X293 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X295 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X297 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X298 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X300 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X305 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X311 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X313 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X314 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X320 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X321 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X325 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X329 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X332 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X335 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X342 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X344 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X345 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X346 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X349 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X351 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X352 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X353 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X356 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X357 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X359 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X365 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X366 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X367 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X368 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X373 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X377 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X383 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X387 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X388 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X389 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X390 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X395 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X398 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X399 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X403 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X406 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X407 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X408 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X410 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X411 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X415 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X422 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X423 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X424 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X425 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X427 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X432 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X435 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X436 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X438 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X440 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X441 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X442 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X443 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X445 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X446 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X448 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X451 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X453 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X455 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X459 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X460 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X466 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X467 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X468 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X470 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X474 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X481 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X483 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X490 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X494 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X501 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X502 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X509 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X511 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X512 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X513 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X514 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X516 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X517 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X521 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X522 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X526 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X528 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X529 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X530 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X532 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X535 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X537 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X538 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X539 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X540 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X544 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X545 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X547 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X548 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X549 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X551 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X552 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X553 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X554 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X555 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X556 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X557 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X562 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X564 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X566 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X569 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X572 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X574 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X577 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X579 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X582 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X583 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X585 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X587 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X588 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X594 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X596 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X598 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X600 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X601 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X602 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X607 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X609 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X610 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X612 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X614 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X619 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X620 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X621 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X622 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X623 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X625 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X626 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X627 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X628 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X630 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X631 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X633 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X634 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X636 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X637 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X639 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X641 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X644 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X646 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33125 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X647 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X650 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X652 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X656 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X661 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X664 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X665 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X668 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X670 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X673 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X674 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X675 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X676 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X678 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X680 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X681 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X683 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X685 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X686 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X688 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X690 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X692 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X693 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X694 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X695 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X696 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X697 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X700 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X701 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X702 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X704 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X705 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X706 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X709 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X713 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X714 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X715 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X717 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X718 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X719 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X720 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X721 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X722 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X725 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X728 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X731 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X736 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X737 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X741 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X743 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X745 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X747 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X748 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X753 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X754 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X755 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X757 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X759 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X760 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X761 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X763 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X764 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X770 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X772 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X773 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X774 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X776 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X778 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X783 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X784 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X786 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X787 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X788 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X790 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X791 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X792 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X793 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X794 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X799 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X801 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X802 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X805 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X806 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X807 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X809 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X810 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X812 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X815 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X816 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X817 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X820 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X823 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X824 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X825 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X827 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X828 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X830 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X831 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X834 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X836 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X839 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X841 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X845 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X846 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X848 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X849 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X851 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X852 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X853 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X854 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X856 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X857 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X858 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X859 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X860 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X861 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X862 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X864 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X868 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X870 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X871 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X878 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X879 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X881 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X882 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X883 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X884 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X885 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X886 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X887 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X888 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X889 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X890 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X892 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X894 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X898 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X899 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X903 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X908 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X912 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X915 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X919 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X921 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X928 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X930 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X932 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X935 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X936 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X941 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X942 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X943 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X946 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X951 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X953 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X954 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X956 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X957 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X958 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X960 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X961 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X965 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X966 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X967 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X968 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X970 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X971 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X972 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X974 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X975 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X977 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X978 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X979 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X984 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X986 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X987 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X989 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X990 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X995 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X997 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X998 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1000 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1001 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1004 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1005 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1007 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1008 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1011 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1014 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1018 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1021 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1022 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1024 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1026 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1030 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1031 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1032 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1034 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1035 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1036 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1037 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1040 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1044 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1045 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1046 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1047 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1048 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1049 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1050 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1053 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1054 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1056 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1057 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1058 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1059 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1061 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1062 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1066 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1068 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1069 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1070 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1071 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1072 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1073 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1075 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1076 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1077 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1081 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1085 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1089 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1091 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1093 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1095 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1096 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1097 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1098 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1100 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1101 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1103 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1104 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1111 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1114 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1115 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1116 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1125 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1128 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1130 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1131 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1132 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1133 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1137 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1141 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1143 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1145 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1146 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1147 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1150 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1153 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1154 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1155 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1158 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1159 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1161 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1162 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1165 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1166 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1173 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1176 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1179 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1182 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1185 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1190 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1193 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1205 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1214 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1215 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1217 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1219 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1222 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1225 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1226 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1231 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1232 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1237 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1243 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1245 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1250 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1259 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1262 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1263 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1266 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1267 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1269 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1270 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1271 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1272 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1277 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1282 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1288 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1291 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1292 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1295 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1315 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1316 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1327 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1329 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1330 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1331 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1332 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1335 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1339 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1343 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1351 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1354 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1358 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1360 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1361 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1365 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1370 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1371 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1372 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1374 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1376 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1378 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1386 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1389 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1392 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1393 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1394 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1395 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1403 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1405 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1408 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1409 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1413 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1416 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1418 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1419 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1426 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1431 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1445 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1460 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1462 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1463 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1464 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1465 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1467 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1469 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1470 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1475 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1476 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1479 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1480 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1483 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1493 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1496 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1497 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1499 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1500 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1504 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1512 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1515 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1516 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1517 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1521 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1528 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1529 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1530 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1532 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1533 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1536 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1538 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1540 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1543 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1544 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1545 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1547 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1548 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1551 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1552 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1553 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1554 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1556 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1557 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1560 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1562 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1567 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1570 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1571 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1572 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1573 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1574 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1577 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1582 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1583 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1585 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1587 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1588 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1589 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1594 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1595 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1598 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1600 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1601 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1602 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1604 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1606 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1610 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1612 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1614 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1617 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1619 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1620 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1621 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1623 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1625 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1626 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1627 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1628 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1630 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1631 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1633 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1634 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1637 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1638 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1639 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1641 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1644 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1645 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1646 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1647 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1649 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1652 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1654 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1656 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1658 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1664 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1665 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1668 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1670 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1673 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1674 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1675 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1676 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1678 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1679 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1680 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1681 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1683 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1685 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1686 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1688 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1690 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1693 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1694 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1695 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1697 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1701 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1702 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1704 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1706 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1707 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1709 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1710 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1713 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1715 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1717 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1718 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1719 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1720 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1721 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1722 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1725 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1727 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1728 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1731 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1733 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1737 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1740 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1741 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1743 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1746 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1747 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1748 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1749 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1751 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1752 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1753 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1754 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1756 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1757 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1761 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1762 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1763 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1765 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1768 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1770 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1772 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1773 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1774 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1777 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1779 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1781 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1783 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1786 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1787 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1788 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1790 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1792 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1793 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1794 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1795 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1799 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1801 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1802 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1803 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1805 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1806 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1807 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1809 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1810 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1812 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1814 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1815 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1817 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1818 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1820 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1821 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1822 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1823 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1824 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1825 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1830 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1831 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1833 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1836 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1838 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1839 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1841 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1844 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1845 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1846 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1847 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1848 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1849 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1850 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1851 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1853 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1854 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1858 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1859 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1860 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1861 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1862 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1864 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1865 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1867 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1868 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1870 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1871 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1872 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1876 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1878 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1882 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1883 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1884 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1886 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1889 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1890 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1892 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1893 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1895 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1899 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1900 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1901 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1903 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1904 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1906 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1908 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1915 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1917 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1919 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1921 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1922 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1932 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1935 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1938 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1941 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1942 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1946 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1948 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1949 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1950 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1954 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1955 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1956 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1958 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1960 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1961 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1965 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1966 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1967 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1968 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1970 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1971 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1972 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1975 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1977 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1978 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1979 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1980 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.33125 ps=9.38 w=4.38 l=0.5
X1981 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1982 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1983 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1984 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1987 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1988 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1989 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1990 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1995 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1996 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1997 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2000 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2001 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2005 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2008 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2011 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2014 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2015 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2016 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2018 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2021 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2022 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2024 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2026 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2027 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2030 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2032 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2034 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2037 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2039 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2040 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2041 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2045 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2046 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2047 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2048 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2053 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2054 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2055 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2056 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2057 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2058 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2059 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2061 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2062 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2063 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2069 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2070 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2071 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2072 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2073 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2074 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2075 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2076 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2077 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2081 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2086 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2087 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2088 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2089 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2091 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2093 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2095 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2096 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2097 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2098 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2109 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2111 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2122 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2124 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2130 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2132 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2139 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2140 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2144 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2153 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2156 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2157 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2165 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2166 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2169 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2178 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2180 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2184 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2185 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2191 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2194 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2195 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2197 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2200 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2205 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2208 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2209 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2217 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2219 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2220 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2221 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2226 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2227 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2228 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2236 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2238 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2239 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2241 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2246 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2248 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2251 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2252 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2254 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2257 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2258 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2260 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2262 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2264 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2265 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2267 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2276 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2278 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2279 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2281 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2286 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2287 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2289 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2296 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2306 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2308 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2318 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2320 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2321 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2322 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2324 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2325 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2330 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2334 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2337 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2339 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2340 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2341 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2347 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2351 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2352 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2353 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2356 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2362 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2363 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2364 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2368 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2369 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2375 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2378 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2386 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2391 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33125 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X2393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2402 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2404 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2406 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2410 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2414 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2421 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2424 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2430 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2434 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2438 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2440 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2444 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2446 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2447 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2450 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2451 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2457 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2458 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2459 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2468 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2472 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2473 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2486 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2487 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2488 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2489 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2490 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2492 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2493 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2499 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2504 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2507 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2509 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2511 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2512 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2516 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2517 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2519 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2521 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2527 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2528 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2529 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2530 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2531 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2532 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2534 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2538 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2540 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2542 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2544 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2545 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2546 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2547 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2548 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2551 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2552 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2553 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2554 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2556 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2557 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2561 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2562 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2563 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2565 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2572 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2574 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2575 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2577 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2578 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2581 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2582 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2583 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2585 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2586 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2587 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2588 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2591 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2592 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2594 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2598 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2599 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2600 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2601 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2602 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2605 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2610 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2611 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2612 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2614 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2619 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2620 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2621 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2623 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2625 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2626 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2627 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2628 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2630 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2631 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2632 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2633 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2634 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2637 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2639 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2641 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2644 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2646 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2647 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2652 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2653 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2656 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2657 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2659 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2663 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2664 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2665 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2668 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2669 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2670 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2672 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2673 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2674 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2675 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2676 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2678 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2680 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2681 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2682 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2683 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2684 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2685 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2686 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2688 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2689 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2690 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2693 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2694 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2695 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2697 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2699 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2701 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2702 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2704 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2706 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2709 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2711 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2712 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2713 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2715 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2717 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2718 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2719 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2720 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2721 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2722 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2725 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2728 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2731 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2737 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2741 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2743 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2747 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2748 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2753 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2754 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2757 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2758 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2761 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2763 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2769 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2770 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2772 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2773 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2774 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2775 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2783 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2786 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2787 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2788 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2789 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2790 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2792 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2793 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2794 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2797 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2799 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2801 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2802 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2805 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2806 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2807 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2809 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2810 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2812 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2815 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2817 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2819 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2820 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2823 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2824 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2825 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2829 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2830 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2831 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2836 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2839 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2841 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2842 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2843 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2845 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2846 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2848 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2849 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2851 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2853 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2854 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2855 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2858 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2859 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2860 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2861 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2862 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2863 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2864 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2868 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2870 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2871 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2878 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2882 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2883 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2884 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2886 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2889 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2890 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2891 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2892 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2897 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2899 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2903 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2905 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2908 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2909 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2910 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2915 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2916 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2919 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2921 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2923 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2932 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2935 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2939 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2941 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2942 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.33125 ps=9.38 w=4.38 l=0.5
X2944 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2946 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2947 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2954 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2956 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2958 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2960 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2961 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2965 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2966 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2967 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2968 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2970 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2971 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2972 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2973 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2975 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2977 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2978 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2979 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2984 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2985 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2987 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2989 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2990 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2995 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2997 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2999 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3000 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3001 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3003 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3005 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3008 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3011 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3012 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3013 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3014 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3018 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3021 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3022 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3023 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3024 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3026 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3028 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3030 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3032 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3034 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3037 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3040 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3042 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3045 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3046 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3047 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3048 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X3051 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3052 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3053 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3054 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3056 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3057 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3058 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3059 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3061 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3062 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3065 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3067 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3069 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3070 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3071 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3072 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3073 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3075 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3076 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3077 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3078 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3079 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3081 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3089 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3091 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3093 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3095 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3096 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3097 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3098 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3106 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3109 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3112 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3114 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3118 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3120 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3121 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3122 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3123 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3126 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3129 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3131 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3133 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3134 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3135 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3137 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3138 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3139 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3140 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3142 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3144 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3148 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3149 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3154 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3159 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3163 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3168 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3175 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3176 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3177 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3178 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3179 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3181 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3186 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3189 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3190 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3192 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3194 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3195 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3196 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3198 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3199 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3201 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3202 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3203 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3210 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3211 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3212 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3215 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3218 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3221 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3227 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3228 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3229 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3230 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3233 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3234 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3243 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3244 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3246 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3247 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3248 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3249 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3250 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3252 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3255 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3256 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3260 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3265 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3269 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3275 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3284 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3289 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3290 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3293 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3294 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3296 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3299 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3300 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3301 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3303 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3306 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3308 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3309 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3310 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3317 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3328 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3333 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3334 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3336 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3337 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3343 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3345 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3350 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3351 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3354 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3360 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3362 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3363 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3364 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3367 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3369 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3370 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3371 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3375 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3376 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3377 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3381 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3384 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3385 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3393 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3394 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3396 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3400 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3402 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3405 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3414 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3415 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3417 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3421 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3425 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3427 a_112_1150# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X3428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3429 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3431 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3432 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3434 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3441 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3442 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3447 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3448 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3452 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3453 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3458 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3461 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3466 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3471 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3474 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3477 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3478 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3480 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3481 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3482 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3484 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3485 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3486 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3487 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3489 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3494 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3496 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3503 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3505 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3506 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3508 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3510 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3512 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3516 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3517 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3518 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3521 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3523 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3524 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3525 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3528 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3529 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3530 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3532 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3538 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3540 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3541 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3544 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3545 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3547 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3548 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3551 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3552 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3553 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3554 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3556 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3557 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3558 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3559 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3562 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3572 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3574 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3576 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3577 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3582 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3583 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3584 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3585 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3587 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3588 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3594 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3597 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3598 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3600 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3601 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3602 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3603 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3608 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3610 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3612 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3613 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3614 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3616 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3619 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3620 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3621 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3623 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3624 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3625 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3626 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3627 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3628 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3630 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3631 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3633 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3634 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3635 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3637 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3639 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3640 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3641 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3642 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3644 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3646 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3647 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3652 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3655 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3656 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3660 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3664 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3665 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3666 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3668 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3670 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3673 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3674 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3675 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3676 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3678 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3680 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3681 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3683 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3685 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3686 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3688 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3690 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3693 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3694 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3695 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3697 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3701 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3702 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3704 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3706 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3708 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3709 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3713 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3715 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3717 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3718 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3719 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3720 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3721 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3722 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3725 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3728 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3729 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3731 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3737 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3738 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3739 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3741 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3742 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3743 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3747 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3748 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3753 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3754 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3757 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3761 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3763 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3770 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3771 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3772 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3773 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3774 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3783 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3785 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3786 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3787 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3788 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3790 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3792 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3793 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3794 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3799 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3800 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3801 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3802 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3804 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3805 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3806 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3807 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3809 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3810 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3812 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3815 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3817 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3820 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3823 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3824 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3825 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3826 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3830 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3831 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3835 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3836 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3837 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3839 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3841 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3845 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3846 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3848 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3849 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3851 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3853 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3854 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3858 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3859 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3860 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3861 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3862 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3864 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3866 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3868 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3869 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3870 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3871 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3873 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3878 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3882 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3883 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3884 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3886 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3889 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3890 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3892 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3899 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3903 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3908 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3914 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3915 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3918 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3919 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3921 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3926 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3927 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3931 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3932 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3934 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3935 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3940 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3941 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3942 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3945 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3946 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3952 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3954 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3956 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3958 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3959 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3960 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3961 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3962 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3964 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3965 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3966 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3967 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3968 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3970 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3971 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3972 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3975 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3977 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3978 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3979 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3984 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3987 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3989 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3990 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3994 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3995 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3997 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4000 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4001 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4005 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4008 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4009 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4010 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4011 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4014 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4017 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4018 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4020 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4021 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4022 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4024 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4026 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4030 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4032 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4034 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4037 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4038 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4040 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4045 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4046 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4047 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4048 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4053 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4054 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4056 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4057 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4058 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4059 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4060 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4061 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4062 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4064 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4069 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4070 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4071 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4072 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4073 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4075 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4076 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4077 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4081 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4082 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4083 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4084 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4089 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4090 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4091 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4093 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4095 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4096 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4097 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4098 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4103 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4105 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4106 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4107 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4113 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4117 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4119 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4125 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4126 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4127 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4128 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4129 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4138 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4142 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4143 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4147 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4150 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4155 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4156 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4158 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4167 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4169 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4170 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4174 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4175 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4177 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4180 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4181 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4187 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4189 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4191 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4199 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4200 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4201 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4202 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4207 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4208 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4209 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4210 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4211 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4212 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4216 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4222 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4224 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4229 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4231 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4235 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4237 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4239 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4240 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4241 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4251 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4254 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4259 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4271 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4274 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4286 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4290 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4291 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4292 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4294 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4298 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4299 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4303 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4307 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4310 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4311 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4312 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4314 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4315 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4316 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4324 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4326 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4327 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4328 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4336 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4340 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4341 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4342 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4344 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4347 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4348 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4349 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4351 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4355 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4361 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4373 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4374 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4379 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4380 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4381 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4382 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4383 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4384 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4387 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4397 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4401 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4404 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4411 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4412 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4413 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4419 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4420 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4422 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4426 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4436 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4437 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4439 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4443 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4444 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4454 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4455 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4457 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4461 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4462 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4463 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4471 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4476 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4479 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4482 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4484 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4485 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4488 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4492 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4495 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4503 a_112_1150# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X4504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4507 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4510 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
.ends

.subckt power_stage p_in sw_node vdd_pwr sky130_fd_sc_hd__inv_4_1/VPB vss dvss
Xsky130_fd_sc_hd__decap_3_0 dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1 dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__inv_4_0 p_in dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ gate_drive_0/in_m sky130_fd_sc_hd__inv_4
Xgate_drive_0 gate_drive_0/in_m gate_drive_0/in_p gate_drive_0/out vdd_pwr vss dvss
+ gate_drive
Xsky130_fd_sc_hd__inv_4_1 gate_drive_0/in_m dvss dvss sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__inv_4_1/VPB gate_drive_0/in_p sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__diode_2_0 p_in dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__diode_2
Xpmos_waffle_48x48_0 vdd_pwr vss gate_drive_0/out sw_node sw_node pmos_waffle_48x48
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RK a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_QRKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_05v0_nvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_nstack itail ena nbias avss vcasc
XXM12 avss avss nbias m1_3726_n2502# sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RK
XXM6 avss vcasc nbias m1_3726_n2502# sky130_fd_pr__nfet_05v0_nvt_QRKT8P
XXM7 avss vcasc ena itail sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__res_high_po_0p35_P35QVK a_380_2984# a_5692_n3416# a_n3770_2984#
+ a_3866_2984# a_3202_n3416# a_n1446_n3416# a_n284_n3416# a_n616_2984# a_4696_n3416#
+ a_4198_2984# a_2206_n3416# a_n1114_2984# a_n4102_2984# a_n616_n3416# a_6190_n3416#
+ a_n6592_2984# a_2372_2984# a_n5762_n3416# a_5360_2984# a_214_2984# a_n3604_2984#
+ a_1210_n3416# a_5194_n3416# a_6522_n3416# a_n4766_n3416# a_1874_2984# a_4862_2984#
+ a_4198_n3416# a_5526_n3416# a_5194_2984# a_n6260_n3416# a_878_n3416# a_n3438_2984#
+ a_n2110_2984# a_n6426_2984# a_2206_2984# a_n118_n3416# a_n3770_n3416# a_4696_2984#
+ a_n5264_n3416# a_48_2984# a_4530_n3416# a_n2774_n3416# a_n1612_2984# a_n4600_2984#
+ a_n5928_2984# a_1708_2984# a_6024_n3416# a_n4268_n3416# a_2870_2984# a_3534_n3416#
+ a_712_2984# a_n1778_n3416# a_5028_2984# a_5028_n3416# a_n948_2984# a_2538_n3416#
+ a_6190_2984# a_n1446_2984# a_n3272_n3416# a_n4434_2984# a_n4600_n3416# a_3202_2984#
+ a_n948_n3416# a_5692_2984# a_380_n3416# a_546_2984# a_4032_n3416# a_n2276_n3416#
+ a_n3604_n3416# a_n3936_2984# a_1542_n3416# a_2704_2984# a_3036_n3416# a_712_n3416#
+ a_n2608_n3416# a_n4268_2984# a_3036_2984# a_6024_2984# a_5858_n3416# a_n1280_n3416#
+ a_n6592_n3416# a_n2442_2984# a_n4102_n3416# a_2538_2984# a_n5430_2984# a_2040_n3416#
+ a_5526_2984# a_1210_2984# a_n1612_n3416# a_n5596_n3416# a_4862_n3416# a_n450_n3416#
+ a_n1944_2984# a_n3106_n3416# a_n4932_2984# a_1044_n3416# a_n450_2984# a_3700_2984#
+ a_6356_n3416# a_214_n3416# a_n5928_n3416# a_n6722_n3546# a_3866_n3416# a_n2276_2984#
+ a_n5264_2984# a_1044_2984# a_4032_2984# a_n2110_n3416# a_n6094_n3416# a_n1778_2984#
+ a_n4766_2984# a_5360_n3416# a_n284_2984# a_3534_2984# a_n4932_n3416# a_6522_2984#
+ a_n1114_n3416# a_2870_n3416# a_n5098_n3416# a_n6426_n3416# a_878_2984# a_4364_n3416#
+ a_n5098_2984# a_n3936_n3416# a_n2940_2984# a_1874_n3416# a_3368_n3416# a_n3272_2984#
+ a_3368_2984# a_48_n3416# a_n6260_2984# a_2040_2984# a_6356_2984# a_n5430_n3416#
+ a_n2940_n3416# a_n118_2984# a_n2774_2984# a_n4434_n3416# a_n5762_2984# a_1542_2984#
+ a_2372_n3416# a_4530_2984# a_5858_2984# a_3700_n3416# a_n1944_n3416# a_n3438_n3416#
+ a_n6094_2984# a_n782_n3416# a_1376_n3416# a_n782_2984# a_2704_n3416# a_546_n3416#
+ a_n3106_2984# a_n1280_2984# a_n5596_2984# a_1376_2984# a_1708_n3416# a_4364_2984#
+ a_n2442_n3416# a_n2608_2984#
X0 a_n3936_2984# a_n3936_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_n1612_2984# a_n1612_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_n6592_2984# a_n6592_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_n4434_2984# a_n4434_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_48_2984# a_48_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_2704_2984# a_2704_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_4862_2984# a_4862_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_3202_2984# a_3202_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_5360_2984# a_5360_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_5526_2984# a_5526_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_n948_2984# a_n948_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_n782_2984# a_n782_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_6024_2984# a_6024_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_n4932_2984# a_n4932_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_1376_2984# a_1376_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_878_2984# a_878_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_4198_2984# a_4198_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_n3770_2984# a_n3770_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_n1446_2984# a_n1446_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_3700_2984# a_3700_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n4268_2984# a_n4268_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n2110_2984# a_n2110_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_1874_2984# a_1874_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_6522_2984# a_6522_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_2372_2984# a_2372_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_2538_2984# a_2538_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_4696_2984# a_4696_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_3036_2984# a_3036_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_5194_2984# a_5194_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_n1944_2984# a_n1944_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_n4766_2984# a_n4766_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n2608_2984# a_n2608_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n2442_2984# a_n2442_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_214_2984# a_214_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n5430_2984# a_n5430_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_n5264_2984# a_n5264_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_n3106_2984# a_n3106_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_2870_2984# a_2870_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_n1280_2984# a_n1280_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_1210_2984# a_1210_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_3534_2984# a_3534_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_5692_2984# a_5692_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_5858_2984# a_5858_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_712_2984# a_712_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_4032_2984# a_4032_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_6190_2984# a_6190_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_6356_2984# a_6356_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_n5928_2984# a_n5928_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_n5762_2984# a_n5762_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n3604_2984# a_n3604_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_n118_2984# a_n118_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_n6426_2984# a_n6426_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_n4102_2984# a_n4102_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_n1778_2984# a_n1778_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_4530_2984# a_4530_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_n4600_2984# a_n4600_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_n2276_2984# a_n2276_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_n5098_2984# a_n5098_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_n616_2984# a_n616_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_1044_2984# a_1044_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_3368_2984# a_3368_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_546_2984# a_546_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_n2940_2984# a_n2940_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_n2774_2984# a_n2774_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_380_2984# a_380_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n5596_2984# a_n5596_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_n3438_2984# a_n3438_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X67 a_n3272_2984# a_n3272_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X68 a_n1114_2984# a_n1114_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X69 a_n6260_2984# a_n6260_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X70 a_n6094_2984# a_n6094_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X71 a_1708_2984# a_1708_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X72 a_1542_2984# a_1542_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X73 a_2206_2984# a_2206_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X74 a_3866_2984# a_3866_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X75 a_2040_2984# a_2040_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X76 a_4364_2984# a_4364_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X77 a_5028_2984# a_5028_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X78 a_n450_2984# a_n450_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X79 a_n284_2984# a_n284_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VPB VPWR X VPWR_uq0 VGND_uq0 VNB
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X4 VGND_uq0 A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR_uq0 a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_772_151# a_404_1133# VGND_uq0 VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X10 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X11 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 VGND_uq0 a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND_uq0 a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_H75TTW a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_pstack pcasc enb itail vcasc pbias avss avdd
XXM13 m1_2150_n1558# avdd pcasc vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__pfet_g5v0d10v5_G8LMTZ_0 itail avdd enb vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss enb sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__pfet_g5v0d10v5_H75TTW_0 m1_2150_n1558# avdd pbias avdd sky130_fd_pr__pfet_g5v0d10v5_H75TTW
.ends

.subckt sky130_fd_pr__res_high_po_0p35_L4QTBM a_3451_2984# a_4447_n3416# a_795_2984#
+ a_1957_n3416# a_n5181_n3416# a_n201_2984# a_n2691_n3416# a_2953_2984# a_n2027_2984#
+ a_n4185_n3416# a_n5015_2984# a_n5513_n3416# a_3451_n3416# a_n1695_n3416# a_3285_2984#
+ a_n3189_n3416# a_n1529_2984# a_n4517_n3416# a_n4517_2984# a_2455_n3416# a_297_n3416#
+ a_n2691_2984# a_2787_2984# a_629_2984# a_n35_2984# a_n865_n3416# a_1459_n3416# a_629_n3416#
+ a_n2193_n3416# a_n3521_n3416# a_n3023_2984# a_n5015_n3416# a_3119_2984# a_n1197_n3416#
+ a_n2525_n3416# a_1293_2984# a_4281_2984# a_n4019_n3416# a_n2525_2984# a_n5513_2984#
+ a_n1529_n3416# a_3783_2984# a_4779_n3416# a_n367_n3416# a_n533_2984# a_n3023_n3416#
+ a_n2359_2984# a_131_n3416# a_n1031_2984# a_n5347_2984# a_1127_2984# a_4115_2984#
+ a_n2027_n3416# a_3783_n3416# a_5277_n3416# a_131_2984# a_n4849_n3416# a_n4849_2984#
+ a_n367_2984# a_n3521_2984# a_n5643_n3546# a_2787_n3416# a_3617_2984# a_1791_2984#
+ a_n1031_n3416# a_4281_n3416# a_n3853_n3416# a_1791_n3416# a_n3355_2984# a_n5347_n3416#
+ a_961_n3416# a_2123_2984# a_3285_n3416# a_4613_n3416# a_5111_2984# a_n201_n3416#
+ a_n2857_n3416# a_n2857_2984# a_2289_n3416# a_1625_2984# a_3617_n3416# a_4613_2984#
+ a_n4351_n3416# a_n699_n3416# a_n3189_2984# a_n1861_n3416# a_n865_2984# a_5111_n3416#
+ a_n3355_n3416# a_1293_n3416# a_2621_n3416# a_n1363_2984# a_n4351_2984# a_463_n3416#
+ a_1459_2984# a_4115_n3416# a_4447_2984# a_n2359_n3416# a_463_2984# a_1625_n3416#
+ a_n699_2984# a_n3853_2984# a_3119_n3416# a_3949_2984# a_2621_2984# a_n1197_2984#
+ a_n1363_n3416# a_n4185_2984# a_297_2984# a_2123_n3416# a_n3687_2984# a_2455_2984#
+ a_5443_2984# a_n533_n3416# a_4945_n3416# a_1127_n3416# a_n1861_2984# a_1957_2984#
+ a_3949_n3416# a_4945_2984# a_n35_n3416# a_n4019_2984# a_n4683_n3416# a_961_2984#
+ a_n2193_2984# a_2289_2984# a_n5181_2984# a_5277_2984# a_5443_n3416# a_n3687_n3416#
+ a_2953_n3416# a_n1695_2984# a_n4683_2984# a_795_n3416# a_4779_2984#
X0 a_n1197_2984# a_n1197_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_3451_2984# a_3451_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_3617_2984# a_3617_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_4115_2984# a_4115_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_2289_2984# a_2289_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_n3521_2984# a_n3521_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_n1695_2984# a_n1695_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_4613_2984# a_4613_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_n2359_2984# a_n2359_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_n2193_2984# a_n2193_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_5111_2984# a_5111_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_n533_2984# a_n533_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_2787_2984# a_2787_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_1127_2984# a_1127_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_3285_2984# a_3285_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_629_2984# a_629_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_n2857_2984# a_n2857_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_n2691_2984# a_n2691_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_463_2984# a_463_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_n3355_2984# a_n3355_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n1031_2984# a_n1031_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n4019_2984# a_n4019_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_n35_2984# a_n35_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_1625_2984# a_1625_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_3949_2984# a_3949_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_2123_2984# a_2123_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_3783_2984# a_3783_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_4447_2984# a_4447_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_961_2984# a_961_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_4281_2984# a_4281_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_n367_2984# a_n367_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n4517_2984# a_n4517_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n3853_2984# a_n3853_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_n5015_2984# a_n5015_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n4351_2984# a_n4351_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_297_2984# a_297_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_2621_2984# a_2621_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_4945_2984# a_4945_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_n3189_2984# a_n3189_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_5443_2984# a_5443_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_n865_2984# a_n865_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_1293_2984# a_1293_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_1459_2984# a_1459_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_n5513_2984# a_n5513_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_795_2984# a_795_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_n3687_2984# a_n3687_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_n1529_2984# a_n1529_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_n1363_2984# a_n1363_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_n4185_2984# a_n4185_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n2027_2984# a_n2027_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_1791_2984# a_1791_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_1957_2984# a_1957_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_n201_2984# a_n201_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_2455_2984# a_2455_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_4779_2984# a_4779_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_3119_2984# a_3119_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_5277_2984# a_5277_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_n1861_2984# a_n1861_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_n699_2984# a_n699_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_n4849_2984# a_n4849_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_n4683_2984# a_n4683_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_n2525_2984# a_n2525_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_131_2984# a_131_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_n5347_2984# a_n5347_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_n5181_2984# a_n5181_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n3023_2984# a_n3023_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_2953_2984# a_2953_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_F3TL5C a_100_n200# a_n292_n422# a_n158_n200# a_n100_n288#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n292_n422# sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_56WC32 a_100_n200# a_n158_n200# a_n332_n422#
+ a_n100_n288#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n332_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QSDYAY w_n487_n497# a_29_n297# a_n287_n200# a_n229_n297#
+ a_229_n200# a_n29_n200#
X0 a_n29_n200# a_n229_n297# a_n287_n200# w_n487_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X1 a_229_n200# a_29_n297# a_n29_n200# w_n487_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_V5WCXY a_n287_n200# a_n487_n288# a_229_n200#
+ a_n545_n200# a_29_n288# a_487_n200# a_n29_n200# a_n229_n288# a_287_n288# a_n679_n422#
X0 a_487_n200# a_287_n288# a_229_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n288# a_n287_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_229_n200# a_29_n288# a_n29_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n287_n200# a_n487_n288# a_n545_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt bias_amp nbias ena inp inn out avss avdd
Xsky130_fd_pr__nfet_05v0_nvt_F3TL5C_0 m1_5615_3673# avss m1_7291_3557# ena sky130_fd_pr__nfet_05v0_nvt_F3TL5C
Xsky130_fd_pr__nfet_g5v0d10v5_56WC32_0 m1_7291_3557# avss avss nbias sky130_fd_pr__nfet_g5v0d10v5_56WC32
Xsky130_fd_pr__pfet_g5v0d10v5_QSDYAY_0 avdd m1_6016_4428# m1_6016_4428# m1_6016_4428#
+ out avdd sky130_fd_pr__pfet_g5v0d10v5_QSDYAY
Xsky130_fd_pr__nfet_g5v0d10v5_V5WCXY_0 m1_6016_4428# inp out m1_5615_3673# inn m1_5615_3673#
+ m1_5615_3673# inp inn avss sky130_fd_pr__nfet_g5v0d10v5_V5WCXY
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MQZGVK m3_n686_n2520# c1_n646_n2480#
X0 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X1 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X2 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X3 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt bias_generator_fe snk_test0 src_test0 vbg ref_in dvdd ena_snk_test0 ena_src_test0
+ bias_amp_0/nbias ref_sel_vbg bias_amp_0/out avdd ena bias_pstack_0[9]/pcasc dvss
+ avss
Xbias_nstack_0[0] snk_test0 ena_test0_3v3 bias_amp_0/nbias avss bias_nstack_0[0]/vcasc
+ bias_nstack
Xbias_nstack_0[1] snk_test0 ena_test0_3v3 bias_amp_0/nbias avss bias_nstack_0[1]/vcasc
+ bias_nstack
Xbias_nstack_0[2] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[3] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[4] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[5] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[6] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[7] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[8] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[9] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[10] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[11] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[12] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[13] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[14] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[15] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[16] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[17] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[18] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[19] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[20] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[21] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[22] bias_amp_0/out enb_vbg_3v3 bias_amp_0/nbias avss bias_nstack_0[22]/vcasc
+ bias_nstack
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 avss vbg sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXR2 m1_26761_7166# m1_31907_766# m1_22445_7166# m1_30081_7166# m1_29583_766# m1_24935_766#
+ m1_25931_766# m1_25765_7166# m1_30911_766# m1_30413_7166# m1_28587_766# m1_25101_7166#
+ m1_22113_7166# m1_25599_766# m1_32571_766# m1_19789_7166# m1_28753_7166# m1_20619_766#
+ m1_31741_7166# m1_26429_7166# m1_22777_7166# m1_27591_766# m1_31575_766# bias_nstack_0[9]/itail
+ m1_21615_766# m1_28089_7166# m1_31077_7166# m1_30579_766# m1_31907_766# m1_31409_7166#
+ m1_19955_766# m1_27259_766# m1_22777_7166# m1_24105_7166# m1_19789_7166# m1_28421_7166#
+ m1_26263_766# m1_22611_766# m1_31077_7166# m1_20951_766# m1_26429_7166# m1_30911_766#
+ m1_23607_766# m1_24769_7166# m1_21781_7166# m1_20453_7166# m1_28089_7166# m1_32239_766#
+ m1_21947_766# m1_29085_7166# m1_29915_766# m1_27093_7166# m1_24603_766# m1_31409_7166#
+ m1_31243_766# m1_25433_7166# m1_28919_766# m1_32405_7166# m1_24769_7166# m1_22943_766#
+ m1_21781_7166# m1_21615_766# m1_29417_7166# m1_25267_766# m1_32073_7166# m1_26595_766#
+ m1_26761_7166# m1_30247_766# m1_23939_766# m1_22611_766# m1_22445_7166# bias_pstack_0[9]/pcasc
+ m1_29085_7166# m1_29251_766# m1_26927_766# m1_23607_766# m1_22113_7166# m1_29417_7166#
+ m1_32405_7166# m1_32239_766# m1_24935_766# ref_in m1_23773_7166# m1_22279_766# m1_28753_7166#
+ m1_20785_7166# m1_28255_766# m1_31741_7166# m1_27425_7166# m1_24603_766# m1_20619_766#
+ m1_31243_766# m1_25931_766# m1_24437_7166# m1_23275_766# m1_21449_7166# m1_27259_766#
+ m1_25765_7166# m1_30081_7166# m1_32571_766# m1_26595_766# m1_20287_766# avss m1_30247_766#
+ m1_24105_7166# m1_21117_7166# m1_27425_7166# m1_30413_7166# m1_24271_766# m1_20287_766#
+ m1_24437_7166# m1_21449_7166# m1_31575_766# m1_26097_7166# m1_29749_7166# m1_21283_766#
+ m1_32737_7166# m1_25267_766# m1_29251_766# m1_21283_766# m1_19955_766# m1_27093_7166#
+ m1_30579_766# m1_21117_7166# m1_22279_766# m1_23441_7166# m1_28255_766# m1_29583_766#
+ m1_23109_7166# m1_29749_7166# m1_26263_766# m1_20121_7166# m1_28421_7166# m1_32737_7166#
+ m1_20951_766# m1_23275_766# m1_26097_7166# m1_23441_7166# m1_21947_766# m1_20453_7166#
+ m1_27757_7166# m1_28587_766# m1_30745_7166# m1_32073_7166# m1_29915_766# m1_24271_766#
+ m1_22943_766# m1_20121_7166# m1_25599_766# m1_27591_766# m1_25433_7166# m1_28919_766#
+ m1_26927_766# m1_23109_7166# m1_25101_7166# m1_20785_7166# m1_27757_7166# bias_pstack_0[9]/pcasc
+ m1_30745_7166# m1_23939_766# m1_23773_7166# sky130_fd_pr__res_high_po_0p35_P35QVK
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0] ena_snk_test0 dvdd dvss avdd avdd ena_test0_3v3
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1] ena_src_test0 dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_2/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2] ena dvdd dvss avdd avdd ena_3v3 avdd dvss dvss
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3] ref_sel_vbg dvdd dvss avdd avdd ena_vbg_3v3 avdd
+ dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__inv_2_2 sky130_fd_sc_hvl__inv_2_2/A dvss dvss avdd avdd enb_test0_3v3
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_4 ena_vbg_3v3 dvss dvss avdd avdd enb_vbg_3v3 sky130_fd_sc_hvl__inv_2
Xbias_pstack_0[0] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[0]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[1] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[1]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[2] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[2]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[3] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[3]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[4] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[4]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[5] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[5]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[6] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[6]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[7] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[7]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[8] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[8]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[9] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[9]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[10] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[10]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[11] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[11]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[12] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[12]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[13] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[13]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[14] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[14]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[15] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[15]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[16] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[16]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[17] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[17]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[18] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[18]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[19] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[19]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[20] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[20]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[21] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[21]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[22] bias_pstack_0[9]/pcasc ena_vbg_3v3 bias_amp_0/out bias_pstack_0[22]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xsky130_fd_pr__res_high_po_0p35_L4QTBM_0 m1_17229_7166# m1_18391_766# m1_14573_7166#
+ m1_15735_766# m1_8763_766# m1_13577_7166# m1_11087_766# m1_16897_7166# m1_11917_7166#
+ m1_9759_766# m1_8929_7166# m1_8431_766# m1_17395_766# m1_12083_766# m1_17229_7166#
+ m1_10755_766# m1_12249_7166# m1_9427_766# m1_9261_7166# m1_16399_766# m1_14075_766#
+ m1_11253_7166# m1_16565_7166# m1_14573_7166# m1_13909_7166# m1_13079_766# m1_15403_766#
+ m1_14407_766# m1_11751_766# m1_10423_766# m1_10921_7166# m1_8763_766# m1_16897_7166#
+ m1_12747_766# m1_11419_766# m1_15237_7166# m1_18225_7166# m1_9759_766# m1_11253_7166#
+ bias_amp_0/inp m1_12415_766# m1_17561_7166# m1_18723_766# m1_13411_766# m1_13245_7166#
+ m1_10755_766# m1_11585_7166# m1_14075_766# m1_12913_7166# m1_8597_7166# m1_14905_7166#
+ m1_17893_7166# m1_11751_766# m1_17727_766# m1_19055_766# m1_13909_7166# m1_9095_766#
+ m1_8929_7166# m1_13577_7166# m1_10257_7166# avss m1_16731_766# m1_17561_7166# m1_15569_7166#
+ m1_12747_766# m1_18059_766# m1_10091_766# m1_15735_766# m1_10589_7166# m1_8431_766#
+ m1_14739_766# m1_15901_7166# m1_17063_766# m1_18391_766# m1_18889_7166# m1_13743_766#
+ m1_11087_766# m1_10921_7166# m1_16067_766# m1_15569_7166# m1_17395_766# m1_18557_7166#
+ m1_9427_766# m1_13079_766# m1_10589_7166# m1_12083_766# m1_12913_7166# m1_19055_766#
+ m1_10423_766# m1_15071_766# m1_16399_766# m1_12581_7166# m1_9593_7166# m1_14407_766#
+ m1_15237_7166# m1_18059_766# m1_18225_7166# m1_11419_766# m1_14241_7166# m1_15403_766#
+ m1_13245_7166# m1_9925_7166# m1_17063_766# m1_17893_7166# m1_16565_7166# m1_12581_7166#
+ m1_12415_766# m1_9593_7166# m1_14241_7166# m1_16067_766# m1_10257_7166# m1_16233_7166#
+ m1_19221_7166# m1_13411_766# m1_18723_766# m1_15071_766# m1_11917_7166# m1_15901_7166#
+ m1_17727_766# m1_18889_7166# m1_13743_766# m1_9925_7166# m1_9095_766# m1_14905_7166#
+ m1_11585_7166# m1_16233_7166# m1_8597_7166# m1_19221_7166# avss m1_10091_766# m1_16731_766#
+ m1_12249_7166# m1_9261_7166# m1_14739_766# m1_18557_7166# sky130_fd_pr__res_high_po_0p35_L4QTBM
Xsky130_fd_sc_hvl__diode_2_0 ena dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_11 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_1 ena_snk_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xbias_amp_0 bias_amp_0/nbias ena_vbg_3v3 bias_amp_0/inp vbg bias_amp_0/out avss avdd
+ bias_amp
Xsky130_fd_sc_hvl__diode_2_2 ena_src_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_3 ref_sel_vbg dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_pr__cap_mim_m3_1_MQZGVK_0 bias_amp_0/inp bias_amp_0/out sky130_fd_pr__cap_mim_m3_1_MQZGVK
Xsky130_fd_pr__cap_mim_m3_1_MQZGVK_1 bias_amp_0/inp bias_amp_0/out sky130_fd_pr__cap_mim_m3_1_MQZGVK
Xsky130_fd_sc_hvl__decap_4_3 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt bias_generator_idac_be avdd dvdd ena[6] ena[3] ena[2] ena[0] ena[1] ena[5]
+ ena[4] ena[7] avss_uq0 avdd_uq0 avdd_uq1 avdd_uq2 a_135144_n10736# m4_89432_13963#
+ a_89514_n1347# m4_89432_n426# a_89514_7744# bias_nstack_3[3]/itail bias_nstack_3[3]/nbias
+ bias_pstack_3[3]/pcasc dvss bias_pstack_2[9]/itail bias_pstack_1[9]/itail bias_pstack_0[9]/itail
+ bias_nstack_1[9]/itail bias_pstack_3[3]/itail bias_nstack_2[9]/itail avss_uq1 bias_nstack_0[9]/itail
+ avss avss_uq2 bias_pstack_3[3]/pbias
Xbias_nstack_0[0] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[0]/vcasc bias_nstack
Xbias_nstack_0[1] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[1]/vcasc bias_nstack
Xbias_nstack_0[2] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[2]/vcasc bias_nstack
Xbias_nstack_0[3] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[3]/vcasc bias_nstack
Xbias_nstack_0[4] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[4]/vcasc bias_nstack
Xbias_nstack_0[5] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[5]/vcasc bias_nstack
Xbias_nstack_0[6] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[6]/vcasc bias_nstack
Xbias_nstack_0[7] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[7]/vcasc bias_nstack
Xbias_nstack_0[8] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[8]/vcasc bias_nstack
Xbias_nstack_0[9] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[9]/vcasc bias_nstack
Xbias_nstack_0[10] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[10]/vcasc bias_nstack
Xbias_nstack_0[11] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[11]/vcasc bias_nstack
Xbias_nstack_0[12] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[12]/vcasc bias_nstack
Xbias_nstack_0[13] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[13]/vcasc bias_nstack
Xbias_nstack_0[14] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[14]/vcasc bias_nstack
Xbias_nstack_0[15] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[15]/vcasc bias_nstack
Xbias_nstack_0[16] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[16]/vcasc bias_nstack
Xbias_nstack_0[17] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[17]/vcasc bias_nstack
Xbias_nstack_0[18] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[18]/vcasc bias_nstack
Xbias_nstack_0[19] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[19]/vcasc bias_nstack
Xbias_nstack_0[20] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[20]/vcasc bias_nstack
Xbias_nstack_0[21] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[21]/vcasc bias_nstack
Xbias_nstack_0[22] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[22]/vcasc bias_nstack
Xbias_nstack_0[23] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[23]/vcasc bias_nstack
Xbias_nstack_0[24] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[24]/vcasc bias_nstack
Xbias_nstack_0[25] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[25]/vcasc bias_nstack
Xbias_nstack_0[26] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[26]/vcasc bias_nstack
Xbias_nstack_0[27] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[27]/vcasc bias_nstack
Xbias_nstack_0[28] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[28]/vcasc bias_nstack
Xbias_nstack_0[29] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[29]/vcasc bias_nstack
Xbias_nstack_0[30] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[30]/vcasc bias_nstack
Xbias_nstack_0[31] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[31]/vcasc bias_nstack
Xbias_nstack_0[32] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[32]/vcasc bias_nstack
Xbias_nstack_0[33] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[33]/vcasc bias_nstack
Xbias_nstack_0[34] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[34]/vcasc bias_nstack
Xbias_nstack_0[35] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[35]/vcasc bias_nstack
Xbias_nstack_0[36] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[36]/vcasc bias_nstack
Xbias_nstack_0[37] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[37]/vcasc bias_nstack
Xbias_nstack_0[38] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[38]/vcasc bias_nstack
Xbias_nstack_0[39] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[39]/vcasc bias_nstack
Xbias_nstack_0[40] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[40]/vcasc bias_nstack
Xbias_nstack_0[41] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[41]/vcasc bias_nstack
Xbias_nstack_0[42] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[42]/vcasc bias_nstack
Xbias_nstack_0[43] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[43]/vcasc bias_nstack
Xbias_nstack_0[44] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[44]/vcasc bias_nstack
Xbias_nstack_0[45] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[45]/vcasc bias_nstack
Xbias_nstack_0[46] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[46]/vcasc bias_nstack
Xbias_nstack_0[47] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[47]/vcasc bias_nstack
Xbias_nstack_0[48] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[48]/vcasc bias_nstack
Xbias_nstack_0[49] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[49]/vcasc bias_nstack
Xbias_nstack_0[50] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[50]/vcasc bias_nstack
Xbias_nstack_0[51] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[51]/vcasc bias_nstack
Xbias_nstack_0[52] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[52]/vcasc bias_nstack
Xbias_nstack_0[53] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[53]/vcasc bias_nstack
Xbias_nstack_0[54] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[54]/vcasc bias_nstack
Xbias_nstack_0[55] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[55]/vcasc bias_nstack
Xbias_nstack_0[56] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[56]/vcasc bias_nstack
Xbias_nstack_0[57] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[57]/vcasc bias_nstack
Xbias_nstack_0[58] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[58]/vcasc bias_nstack
Xbias_nstack_0[59] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[59]/vcasc bias_nstack
Xbias_nstack_0[60] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[60]/vcasc bias_nstack
Xbias_nstack_0[61] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[61]/vcasc bias_nstack
Xbias_nstack_0[62] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[62]/vcasc bias_nstack
Xbias_nstack_0[63] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[63]/vcasc bias_nstack
Xbias_nstack_0[64] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[64]/vcasc bias_nstack
Xbias_nstack_0[65] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[65]/vcasc bias_nstack
Xbias_nstack_0[66] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[66]/vcasc bias_nstack
Xbias_nstack_0[67] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[67]/vcasc bias_nstack
Xbias_nstack_0[68] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[68]/vcasc bias_nstack
Xbias_nstack_0[69] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[69]/vcasc bias_nstack
Xbias_nstack_0[70] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[70]/vcasc bias_nstack
Xbias_nstack_0[71] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[71]/vcasc bias_nstack
Xbias_nstack_0[72] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[72]/vcasc bias_nstack
Xbias_nstack_0[73] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[73]/vcasc bias_nstack
Xbias_nstack_0[74] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[74]/vcasc bias_nstack
Xbias_nstack_0[75] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[75]/vcasc bias_nstack
Xbias_nstack_1[0] bias_nstack_1[9]/itail avss_uq1 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[0]/vcasc bias_nstack
Xbias_nstack_1[1] bias_nstack_1[9]/itail bias_nstack_1[1]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[1]/vcasc bias_nstack
Xbias_nstack_1[2] bias_nstack_1[9]/itail bias_nstack_1[3]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[2]/vcasc bias_nstack
Xbias_nstack_1[3] bias_nstack_1[9]/itail bias_nstack_1[3]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[3]/vcasc bias_nstack
Xbias_nstack_1[4] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[4]/vcasc bias_nstack
Xbias_nstack_1[5] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[5]/vcasc bias_nstack
Xbias_nstack_1[6] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[6]/vcasc bias_nstack
Xbias_nstack_1[7] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[7]/vcasc bias_nstack
Xbias_nstack_1[8] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[8]/vcasc bias_nstack
Xbias_nstack_1[9] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[9]/vcasc bias_nstack
Xbias_nstack_1[10] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[10]/vcasc bias_nstack
Xbias_nstack_1[11] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[11]/vcasc bias_nstack
Xbias_nstack_1[12] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[12]/vcasc bias_nstack
Xbias_nstack_1[13] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[13]/vcasc bias_nstack
Xbias_nstack_1[14] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[14]/vcasc bias_nstack
Xbias_nstack_1[15] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[15]/vcasc bias_nstack
Xbias_nstack_1[16] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[16]/vcasc bias_nstack
Xbias_nstack_1[17] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[17]/vcasc bias_nstack
Xbias_nstack_1[18] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[18]/vcasc bias_nstack
Xbias_nstack_1[19] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[19]/vcasc bias_nstack
Xbias_nstack_1[20] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[20]/vcasc bias_nstack
Xbias_nstack_1[21] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[21]/vcasc bias_nstack
Xbias_nstack_1[22] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[22]/vcasc bias_nstack
Xbias_nstack_1[23] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[23]/vcasc bias_nstack
Xbias_nstack_1[24] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[24]/vcasc bias_nstack
Xbias_nstack_1[25] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[25]/vcasc bias_nstack
Xbias_nstack_1[26] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[26]/vcasc bias_nstack
Xbias_nstack_1[27] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[27]/vcasc bias_nstack
Xbias_nstack_1[28] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[28]/vcasc bias_nstack
Xbias_nstack_1[29] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[29]/vcasc bias_nstack
Xbias_nstack_1[30] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[30]/vcasc bias_nstack
Xbias_nstack_1[31] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[31]/vcasc bias_nstack
Xbias_nstack_1[32] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[32]/vcasc bias_nstack
Xbias_nstack_1[33] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[33]/vcasc bias_nstack
Xbias_nstack_1[34] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[34]/vcasc bias_nstack
Xbias_nstack_1[35] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[35]/vcasc bias_nstack
Xbias_nstack_1[36] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[36]/vcasc bias_nstack
Xbias_nstack_1[37] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[37]/vcasc bias_nstack
Xbias_nstack_1[38] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[38]/vcasc bias_nstack
Xbias_nstack_1[39] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[39]/vcasc bias_nstack
Xbias_nstack_1[40] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[40]/vcasc bias_nstack
Xbias_nstack_1[41] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[41]/vcasc bias_nstack
Xbias_nstack_1[42] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[42]/vcasc bias_nstack
Xbias_nstack_1[43] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[43]/vcasc bias_nstack
Xbias_nstack_1[44] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[44]/vcasc bias_nstack
Xbias_nstack_1[45] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[45]/vcasc bias_nstack
Xbias_nstack_1[46] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[46]/vcasc bias_nstack
Xbias_nstack_1[47] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[47]/vcasc bias_nstack
Xbias_nstack_1[48] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[48]/vcasc bias_nstack
Xbias_nstack_1[49] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[49]/vcasc bias_nstack
Xbias_nstack_1[50] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[50]/vcasc bias_nstack
Xbias_nstack_1[51] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[51]/vcasc bias_nstack
Xbias_nstack_1[52] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[52]/vcasc bias_nstack
Xbias_nstack_1[53] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[53]/vcasc bias_nstack
Xbias_nstack_1[54] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[54]/vcasc bias_nstack
Xbias_nstack_1[55] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[55]/vcasc bias_nstack
Xbias_nstack_1[56] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[56]/vcasc bias_nstack
Xbias_nstack_1[57] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[57]/vcasc bias_nstack
Xbias_nstack_1[58] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[58]/vcasc bias_nstack
Xbias_nstack_1[59] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[59]/vcasc bias_nstack
Xbias_nstack_1[60] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[60]/vcasc bias_nstack
Xbias_nstack_1[61] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[61]/vcasc bias_nstack
Xbias_nstack_1[62] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[62]/vcasc bias_nstack
Xbias_nstack_1[63] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[63]/vcasc bias_nstack
Xbias_nstack_1[64] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[64]/vcasc bias_nstack
Xbias_nstack_1[65] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[65]/vcasc bias_nstack
Xbias_nstack_1[66] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[66]/vcasc bias_nstack
Xbias_nstack_1[67] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[67]/vcasc bias_nstack
Xbias_nstack_1[68] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[68]/vcasc bias_nstack
Xbias_nstack_1[69] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[69]/vcasc bias_nstack
Xbias_nstack_1[70] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[70]/vcasc bias_nstack
Xbias_nstack_1[71] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[71]/vcasc bias_nstack
Xbias_nstack_1[72] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[72]/vcasc bias_nstack
Xbias_nstack_1[73] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[73]/vcasc bias_nstack
Xbias_nstack_1[74] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[74]/vcasc bias_nstack
Xbias_nstack_1[75] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[75]/vcasc bias_nstack
Xbias_nstack_1[76] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[76]/vcasc bias_nstack
Xbias_nstack_1[77] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[77]/vcasc bias_nstack
Xbias_nstack_1[78] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[78]/vcasc bias_nstack
Xbias_nstack_1[79] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[79]/vcasc bias_nstack
Xbias_nstack_1[80] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[80]/vcasc bias_nstack
Xbias_nstack_1[81] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[81]/vcasc bias_nstack
Xbias_nstack_1[82] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[82]/vcasc bias_nstack
Xbias_nstack_1[83] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[83]/vcasc bias_nstack
Xbias_nstack_1[84] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[84]/vcasc bias_nstack
Xbias_nstack_1[85] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[85]/vcasc bias_nstack
Xbias_nstack_1[86] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[86]/vcasc bias_nstack
Xbias_nstack_1[87] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[87]/vcasc bias_nstack
Xsky130_fd_sc_hvl__decap_4_8 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xbias_nstack_2[0] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[0]/vcasc
+ bias_nstack
Xbias_nstack_2[1] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[1]/vcasc
+ bias_nstack
Xbias_nstack_2[2] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[2]/vcasc
+ bias_nstack
Xbias_nstack_2[3] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[3]/vcasc
+ bias_nstack
Xbias_nstack_2[4] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[4]/vcasc
+ bias_nstack
Xbias_nstack_2[5] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[5]/vcasc
+ bias_nstack
Xbias_nstack_2[6] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[6]/vcasc
+ bias_nstack
Xbias_nstack_2[7] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[7]/vcasc
+ bias_nstack
Xbias_nstack_2[8] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[8]/vcasc
+ bias_nstack
Xbias_nstack_2[9] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[9]/vcasc
+ bias_nstack
Xbias_nstack_2[10] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[10]/vcasc
+ bias_nstack
Xbias_nstack_2[11] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[11]/vcasc
+ bias_nstack
Xbias_nstack_2[12] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[12]/vcasc
+ bias_nstack
Xbias_nstack_2[13] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[13]/vcasc
+ bias_nstack
Xbias_nstack_2[14] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[14]/vcasc
+ bias_nstack
Xbias_nstack_2[15] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[15]/vcasc
+ bias_nstack
Xbias_nstack_2[16] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[16]/vcasc
+ bias_nstack
Xbias_nstack_2[17] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[17]/vcasc
+ bias_nstack
Xbias_nstack_2[18] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[18]/vcasc
+ bias_nstack
Xbias_nstack_2[19] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[19]/vcasc
+ bias_nstack
Xbias_nstack_2[20] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[20]/vcasc
+ bias_nstack
Xbias_nstack_2[21] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[21]/vcasc
+ bias_nstack
Xbias_nstack_2[22] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[22]/vcasc
+ bias_nstack
Xbias_nstack_2[23] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[23]/vcasc
+ bias_nstack
Xbias_nstack_2[24] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[24]/vcasc
+ bias_nstack
Xbias_nstack_2[25] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[25]/vcasc
+ bias_nstack
Xbias_nstack_2[26] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[26]/vcasc
+ bias_nstack
Xbias_nstack_2[27] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[27]/vcasc
+ bias_nstack
Xbias_nstack_2[28] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[28]/vcasc
+ bias_nstack
Xbias_nstack_2[29] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[29]/vcasc
+ bias_nstack
Xbias_nstack_2[30] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[30]/vcasc
+ bias_nstack
Xbias_nstack_2[31] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[31]/vcasc
+ bias_nstack
Xbias_nstack_2[32] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[32]/vcasc
+ bias_nstack
Xbias_nstack_2[33] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[33]/vcasc
+ bias_nstack
Xbias_nstack_2[34] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[34]/vcasc
+ bias_nstack
Xbias_nstack_2[35] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[35]/vcasc
+ bias_nstack
Xbias_nstack_2[36] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[36]/vcasc
+ bias_nstack
Xbias_nstack_2[37] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[37]/vcasc
+ bias_nstack
Xbias_nstack_2[38] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[38]/vcasc
+ bias_nstack
Xbias_nstack_2[39] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[39]/vcasc
+ bias_nstack
Xbias_nstack_2[40] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[40]/vcasc
+ bias_nstack
Xbias_nstack_2[41] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[41]/vcasc
+ bias_nstack
Xbias_nstack_2[42] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[42]/vcasc
+ bias_nstack
Xbias_nstack_2[43] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[43]/vcasc
+ bias_nstack
Xbias_nstack_2[44] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[44]/vcasc
+ bias_nstack
Xbias_nstack_2[45] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[45]/vcasc
+ bias_nstack
Xbias_nstack_2[46] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[46]/vcasc
+ bias_nstack
Xbias_nstack_2[47] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[47]/vcasc
+ bias_nstack
Xbias_nstack_2[48] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[48]/vcasc
+ bias_nstack
Xbias_nstack_2[49] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[49]/vcasc
+ bias_nstack
Xbias_nstack_2[50] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[50]/vcasc
+ bias_nstack
Xbias_nstack_2[51] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[51]/vcasc
+ bias_nstack
Xbias_nstack_2[52] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[52]/vcasc
+ bias_nstack
Xbias_nstack_2[53] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[53]/vcasc
+ bias_nstack
Xbias_nstack_2[54] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[54]/vcasc
+ bias_nstack
Xbias_nstack_2[55] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[55]/vcasc
+ bias_nstack
Xbias_nstack_2[56] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[56]/vcasc
+ bias_nstack
Xbias_nstack_2[57] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[57]/vcasc
+ bias_nstack
Xbias_nstack_2[58] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[58]/vcasc
+ bias_nstack
Xbias_nstack_2[59] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[59]/vcasc
+ bias_nstack
Xbias_nstack_2[60] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[60]/vcasc
+ bias_nstack
Xbias_nstack_2[61] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[61]/vcasc
+ bias_nstack
Xbias_nstack_2[62] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[62]/vcasc
+ bias_nstack
Xbias_nstack_2[63] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[63]/vcasc
+ bias_nstack
Xbias_nstack_2[64] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[64]/vcasc
+ bias_nstack
Xbias_nstack_2[65] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[65]/vcasc
+ bias_nstack
Xbias_nstack_2[66] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[66]/vcasc
+ bias_nstack
Xbias_nstack_2[67] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[67]/vcasc
+ bias_nstack
Xbias_nstack_2[68] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[68]/vcasc
+ bias_nstack
Xbias_nstack_2[69] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[69]/vcasc
+ bias_nstack
Xbias_nstack_2[70] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[70]/vcasc
+ bias_nstack
Xbias_nstack_2[71] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[71]/vcasc
+ bias_nstack
Xbias_nstack_2[72] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[72]/vcasc
+ bias_nstack
Xbias_nstack_2[73] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[73]/vcasc
+ bias_nstack
Xbias_nstack_2[74] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[74]/vcasc
+ bias_nstack
Xbias_nstack_2[75] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[75]/vcasc
+ bias_nstack
Xbias_nstack_2[76] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[76]/vcasc
+ bias_nstack
Xbias_nstack_2[77] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[77]/vcasc
+ bias_nstack
Xbias_nstack_2[78] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[78]/vcasc
+ bias_nstack
Xbias_nstack_2[79] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[79]/vcasc
+ bias_nstack
Xbias_nstack_2[80] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[80]/vcasc
+ bias_nstack
Xbias_nstack_2[81] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[81]/vcasc
+ bias_nstack
Xbias_nstack_2[82] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[82]/vcasc
+ bias_nstack
Xbias_nstack_2[83] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[83]/vcasc
+ bias_nstack
Xbias_nstack_2[84] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[84]/vcasc
+ bias_nstack
Xbias_nstack_2[85] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[85]/vcasc
+ bias_nstack
Xbias_nstack_2[86] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[86]/vcasc
+ bias_nstack
Xbias_nstack_2[87] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[87]/vcasc
+ bias_nstack
Xsky130_fd_sc_hvl__decap_4_9 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xbias_nstack_3[0] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[0]/vcasc bias_nstack
Xbias_nstack_3[1] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[1]/vcasc bias_nstack
Xbias_nstack_3[2] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[2]/vcasc bias_nstack
Xbias_nstack_3[3] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[3]/vcasc bias_nstack
Xsky130_fd_sc_hvl__inv_2_0 ena_bit7 dvss dvss avdd_uq2 avdd_uq2 enb_bit7 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 ena_bit3 dvss dvss avdd_uq2 avdd_uq2 enb_bit3 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] ena[7] dvdd dvss avdd_uq2 avdd_uq2 ena_bit7
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] ena[6] dvdd dvss avdd_uq2 avdd_uq2 ena_bit6
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|0] ena[5] dvdd dvss avdd_uq2 avdd_uq2 ena_bit5
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|0] ena[4] dvdd dvss avdd_uq2 avdd_uq2 ena_bit4
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] ena[3] dvdd dvss avdd_uq2 avdd_uq2 ena_bit3
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] ena[2] dvdd dvss avdd_uq2 avdd_uq2 ena_bit2
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|1] ena[1] dvdd dvss avdd_uq2 avdd_uq2 bias_nstack_1[3]/ena
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|1] ena[0] dvdd dvss avdd_uq2 avdd_uq2 bias_nstack_1[1]/ena
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__inv_2_3 ena_bit5 dvss dvss avdd_uq2 avdd_uq2 enb_bit5 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_2 ena_bit6 dvss dvss avdd_uq2 avdd_uq2 enb_bit6 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_4 bias_nstack_1[1]/ena dvss dvss avdd_uq2 avdd_uq2 bias_pstack_1[1]/enb
+ sky130_fd_sc_hvl__inv_2
Xbias_pstack_0[0] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[1] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[1]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[2] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[2]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[3] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[3]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[4] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[4]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[5] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[5]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[6] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[6]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[7] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[7]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[8] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[8]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[9] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[9]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[10] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[10]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[11] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[11]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[12] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[12]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[13] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[13]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[14] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[14]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[15] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[15]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[16] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[16]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[17] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[17]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[18] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[18]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[19] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[19]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[20] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[20]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[21] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[21]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[22] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[22]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[23] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[23]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[24] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[24]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[25] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[25]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[26] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[26]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[27] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[27]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[28] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[28]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[29] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[29]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[30] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[30]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[31] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[31]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[32] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[32]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[33] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[33]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[34] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[34]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[35] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[35]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[36] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[36]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[37] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[37]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[38] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[38]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[39] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[39]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[40] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[40]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[41] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[41]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[42] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[42]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[43] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[43]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[44] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[44]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[45] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[45]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[46] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[46]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[47] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[47]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[48] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[48]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[49] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[49]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[50] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[50]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[51] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[51]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[52] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[52]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[53] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[53]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[54] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[54]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[55] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[55]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[56] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[56]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[57] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[57]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[58] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[58]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[59] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[59]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[60] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[60]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[61] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[61]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[62] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[62]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[63] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[63]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[64] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[64]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[65] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[65]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[66] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[66]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[67] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[67]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[68] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[68]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[69] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[69]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[70] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[70]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[71] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[71]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[72] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[72]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[73] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[73]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[74] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[74]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[75] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[75]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_1[0] bias_pstack_3[3]/pcasc avdd_uq1 bias_pstack_1[9]/itail bias_pstack_1[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[1] bias_pstack_3[3]/pcasc bias_pstack_1[1]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[1]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[2] bias_pstack_3[3]/pcasc bias_pstack_1[3]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[2]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[3] bias_pstack_3[3]/pcasc bias_pstack_1[3]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[3]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[4] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[4]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[5] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[5]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[6] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[6]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[7] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[7]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[8] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[8]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[9] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[9]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[10] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[10]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[11] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[11]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[12] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[12]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[13] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[13]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[14] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[14]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[15] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[15]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[16] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[16]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[17] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[17]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[18] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[18]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[19] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[19]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[20] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[20]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[21] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[21]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[22] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[22]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[23] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[23]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[24] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[24]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[25] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[25]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[26] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[26]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[27] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[27]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[28] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[28]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[29] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[29]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[30] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[30]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[31] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[31]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[32] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[32]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[33] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[33]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[34] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[34]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[35] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[35]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[36] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[36]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[37] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[37]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[38] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[38]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[39] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[39]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[40] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[40]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[41] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[41]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[42] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[42]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[43] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[43]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[44] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[44]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[45] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[45]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[46] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[46]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[47] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[47]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[48] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[48]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[49] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[49]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[50] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[50]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[51] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[51]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[52] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[52]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[53] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[53]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[54] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[54]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[55] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[55]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[56] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[56]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[57] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[57]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[58] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[58]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[59] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[59]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[60] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[60]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[61] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[61]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[62] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[62]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[63] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[63]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[64] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[64]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[65] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[65]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[66] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[66]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[67] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[67]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[68] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[68]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[69] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[69]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[70] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[70]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[71] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[71]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[72] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[72]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[73] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[73]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[74] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[74]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[75] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[75]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[76] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[76]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[77] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[77]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[78] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[78]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[79] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[79]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[80] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[80]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[81] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[81]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[82] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[82]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[83] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[83]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[84] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[84]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[85] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[85]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[86] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[86]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[87] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[87]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_2[0] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[0]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[1] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[1]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[2] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[2]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[3] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[3]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[4] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[4]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[5] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[5]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[6] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[6]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[7] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[7]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[8] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[8]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[9] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[9]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[10] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[10]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[11] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[11]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[12] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[12]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[13] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[13]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[14] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[14]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[15] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[15]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[16] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[16]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[17] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[17]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[18] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[18]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[19] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[19]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[20] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[20]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[21] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[21]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[22] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[22]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[23] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[23]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[24] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[24]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[25] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[25]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[26] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[26]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[27] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[27]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[28] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[28]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[29] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[29]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[30] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[30]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[31] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[31]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[32] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[32]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[33] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[33]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[34] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[34]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[35] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[35]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[36] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[36]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[37] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[37]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[38] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[38]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[39] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[39]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[40] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[40]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[41] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[41]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[42] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[42]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[43] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[43]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[44] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[44]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[45] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[45]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[46] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[46]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[47] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[47]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[48] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[48]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[49] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[49]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[50] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[50]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[51] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[51]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[52] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[52]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[53] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[53]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[54] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[54]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[55] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[55]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[56] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[56]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[57] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[57]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[58] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[58]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[59] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[59]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[60] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[60]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[61] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[61]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[62] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[62]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[63] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[63]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[64] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[64]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[65] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[65]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[66] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[66]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[67] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[67]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[68] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[68]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[69] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[69]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[70] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[70]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[71] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[71]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[72] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[72]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[73] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[73]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[74] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[74]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[75] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[75]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[76] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[76]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[77] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[77]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[78] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[78]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[79] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[79]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[80] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[80]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[81] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[81]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[82] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[82]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[83] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[83]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[84] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[84]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[85] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[85]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[86] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[86]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[87] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[87]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xsky130_fd_sc_hvl__inv_2_7 ena_bit2 dvss dvss avdd_uq2 avdd_uq2 enb_bit2 sky130_fd_sc_hvl__inv_2
Xbias_pstack_3[0] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[1] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[1]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[2] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[2]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[3] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[3]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xsky130_fd_sc_hvl__decap_4_10 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_0 ena[3] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_11 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_1 ena[7] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_13 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_12 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_2 ena[0] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_3 ena[4] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_4 ena[1] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_16 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_5 ena[5] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_17 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_6 ena[2] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_10 ena_bit4 dvss dvss avdd_uq2 avdd_uq2 enb_bit4 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_7 ena[6] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_11 bias_nstack_1[3]/ena dvss dvss avdd_uq2 avdd_uq2 bias_pstack_1[3]/enb
+ sky130_fd_sc_hvl__inv_2
.ends

.subckt sky130_ef_ip__idac3v_8bit din[6] din[3] din[2] din[0] din[1] din[5] din[4]
+ din[7] ref_sel_vbg ena vbg snk_out src_out ref_in avdd dvdd avss dvss
Xbias_generator_fe_0 bias_generator_fe_0/snk_test0 bias_generator_fe_0/src_test0 vbg
+ ref_in dvdd dvss dvss bias_generator_fe_0/bias_amp_0/nbias ref_sel_vbg bias_generator_fe_0/bias_amp_0/out
+ avdd ena bias_generator_fe_0/bias_pstack_0[9]/pcasc dvss avss bias_generator_fe
Xbias_generator_idac_be_0 avdd dvdd din[6] din[3] din[2] din[0] din[1] din[5] din[4]
+ din[7] avss avdd avdd avdd dvss dvdd dvss dvdd dvss snk_out bias_generator_fe_0/bias_amp_0/nbias
+ bias_generator_fe_0/bias_pstack_0[9]/pcasc dvss src_out src_out src_out snk_out
+ src_out snk_out avss snk_out avss avss bias_generator_fe_0/bias_amp_0/out bias_generator_idac_be
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BWAZV5 a_n700_n197# a_700_n100# w_n958_n397#
+ a_n758_n100#
X0 a_700_n100# a_n700_n197# a_n758_n100# w_n958_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_A2FZRM a_n900_n188# a_n900_n1024# a_900_n518#
+ a_n900_648# a_n958_318# a_n958_n518# a_900_736# a_n1102_n1158# a_900_n100# a_900_n936#
+ a_900_318# a_n900_230# a_n958_n100# a_n958_736# a_n958_n936# a_n900_n606#
X0 a_900_n100# a_n900_n188# a_n958_n100# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X1 a_900_n518# a_n900_n606# a_n958_n518# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X2 a_900_318# a_n900_230# a_n958_318# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X3 a_900_n936# a_n900_n1024# a_n958_n936# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X4 a_900_736# a_n900_648# a_n958_736# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6 a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PC2PN5 w_n1258_n397# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1258_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69K6TN a_700_n100# a_n758_n100# a_n700_n188#
+ a_n902_n322#
X0 a_700_n100# a_n700_n188# a_n758_n100# a_n902_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QZEXQH a_1044_n1416# a_214_n1416# a_n1114_n1416#
+ a_546_984# a_n1114_984# a_n118_984# a_48_n1416# a_1376_n1416# a_n450_984# a_n782_n1416#
+ a_878_984# a_546_n1416# a_n1446_984# a_712_984# a_n1446_n1416# a_n284_n1416# a_n616_n1416#
+ a_n782_984# a_1210_n1416# a_1044_984# a_878_n1416# a_n118_n1416# a_n616_984# a_48_984#
+ a_380_984# a_1376_984# a_n948_n1416# a_n1576_n1546# a_380_n1416# a_n948_984# a_712_n1416#
+ a_1210_984# a_214_984# a_n1280_n1416# a_n284_984# a_n450_n1416# a_n1280_984#
X0 a_n1280_984# a_n1280_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n948_984# a_n948_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_1210_984# a_1210_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n616_984# a_n616_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_380_984# a_380_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_878_984# a_878_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_546_984# a_546_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_n1446_984# a_n1446_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_1376_984# a_1376_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_214_984# a_214_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_n1114_984# a_n1114_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n284_984# a_n284_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_1044_984# a_1044_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_n450_984# a_n450_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_48_984# a_48_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_712_984# a_712_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_n782_984# a_n782_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_n118_984# a_n118_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H a_1044_n1416# a_214_n1416# a_n2276_984#
+ a_n2110_n1416# a_1542_984# a_n1114_n1416# a_2870_n1416# a_546_984# a_n1114_984#
+ a_n118_984# a_n2110_984# a_1874_n1416# a_2538_984# a_48_n1416# a_n2940_n1416# a_2372_n1416#
+ a_n1944_n1416# a_1874_984# a_n782_n1416# a_n450_984# a_1376_n1416# a_2870_984# a_878_984#
+ a_2704_n1416# a_546_n1416# a_n1446_984# a_n2442_984# a_1708_n1416# a_n2442_n1416#
+ a_n1446_n1416# a_712_984# a_n284_n1416# a_1708_984# a_2206_n1416# a_2704_984# a_n782_984#
+ a_n616_n1416# a_n1778_984# a_n2774_984# a_1210_n1416# a_1044_984# a_2040_984# a_n1612_984#
+ a_878_n1416# a_n118_n1416# a_n616_984# a_n2774_n1416# a_n2608_984# a_n1778_n1416#
+ a_48_984# a_2538_n1416# a_380_984# a_1376_984# a_n948_n1416# a_2372_984# a_n1944_984#
+ a_380_n1416# a_n2276_n1416# a_n948_984# a_n3070_n1546# a_n2940_984# a_1542_n1416#
+ a_712_n1416# a_n2608_n1416# a_1210_984# a_n1280_n1416# a_214_984# a_2040_n1416#
+ a_n1612_n1416# a_n1280_984# a_2206_984# a_n450_n1416# a_n284_984#
X0 a_1542_984# a_1542_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n1280_984# a_n1280_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_n948_984# a_n948_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_2704_984# a_2704_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_1210_984# a_1210_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_1708_984# a_1708_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_n616_984# a_n616_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_n2774_984# a_n2774_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n2110_984# a_n2110_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_380_984# a_380_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_878_984# a_878_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n1778_984# a_n1778_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_n2442_984# a_n2442_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_n2940_984# a_n2940_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_546_984# a_546_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_n1446_984# a_n1446_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_2372_984# a_2372_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_1376_984# a_1376_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X18 a_n2608_984# a_n2608_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X19 a_214_984# a_214_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X20 a_n1114_984# a_n1114_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X21 a_n284_984# a_n284_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X22 a_2040_984# a_2040_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X23 a_2538_984# a_2538_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X24 a_1044_984# a_1044_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X25 a_n1944_984# a_n1944_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X26 a_n450_984# a_n450_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X27 a_48_984# a_48_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X28 a_2206_984# a_2206_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X29 a_2870_984# a_2870_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X30 a_712_984# a_712_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X31 a_1874_984# a_1874_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X32 a_n1612_984# a_n1612_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X33 a_n782_984# a_n782_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X34 a_n2276_984# a_n2276_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X35 a_n118_984# a_n118_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_743D3R a_n248_n2546# a_48_n2416# a_n118_1984#
+ a_n118_n2416# a_48_1984#
X0 a_48_1984# a_48_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X1 a_n118_1984# a_n118_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MRZGNS c1_n1646_n1500# m3_n1686_n1540#
X0 c1_n1646_n1500# m3_n1686_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S__0 m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PXBJUB a_n1000_n188# a_n1192_n322# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1192_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_47NWVV a_n258_n100# a_n200_n197# a_200_n100#
+ w_n458_n397#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n458_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YHRXVR a_n129_n2415# a_819_2457# a_n977_2545#
+ a_n1609_n4763# a_n1135_n1109# a_n1551_21# a_n503_n4763# a_603_n3545# a_1235_109#
+ a_n1609_n1109# a_n29_4981# a_445_3763# a_n1135_109# a_n1077_2457# a_n1235_n2415#
+ a_n503_n1109# a_1393_4981# a_n29_1327# a_345_2457# a_1235_n3545# a_977_n3633# a_n761_3675#
+ a_n603_n2415# a_1393_1327# a_1293_3675# a_n919_2457# a_977_21# a_n345_n4763# a_445_n3545#
+ a_n503_2545# a_129_2545# a_n1077_n2415# a_n187_4981# a_n1293_2545# a_n819_n4763#
+ a_919_n3545# a_n345_n1109# a_n1551_3675# a_187_21# a_1077_3763# a_n1451_n4763# a_29_n4851#
+ a_1077_n3545# a_977_2457# a_n187_1327# a_n819_n1109# a_503_n2415# a_n129_n1197#
+ a_n445_n2415# a_n445_2457# a_n1451_n1109# a_n977_109# a_1077_109# a_n919_n2415#
+ a_n1235_n1197# a_1135_n2415# a_n1551_n2415# a_29_4893# a_n187_n4763# a_287_n3545#
+ a_1451_21# a_29_1239# a_1551_n3545# a_n187_n1109# a_603_3763# a_n603_n1197# a_n1293_n4763#
+ a_n1235_2457# a_n129_4893# a_345_n2415# a_1551_4981# a_n287_n2415# a_129_109# a_n1293_n1109#
+ a_n129_1239# a_503_2457# a_n661_2545# a_n445_21# a_819_n2415# a_29_n6069# a_287_2545#
+ a_n661_n4763# a_761_n3545# a_1551_1327# a_n819_4981# a_n29_n3545# a_187_4893# a_1451_3675#
+ a_n1077_n1197# a_n1393_n2415# a_n661_n1109# a_n819_1327# a_187_1239# a_1393_n3545#
+ a_503_n1197# a_n445_n1197# a_n761_n2415# a_n345_4981# a_n1451_2545# a_187_n2415#
+ a_n919_n1197# a_n1609_109# a_n1609_4981# a_1235_3763# a_1135_n1197# a_n345_1327#
+ a_n1551_n1197# a_1451_n2415# a_n603_2457# a_n1609_1327# a_129_n5981# a_1135_2457#
+ a_n1077_21# a_761_3763# a_n977_n4763# a_n1393_2457# a_n287_4893# a_129_n2327# a_345_n1197#
+ a_n1135_4981# a_n977_n1109# a_661_n2415# a_n287_1239# a_661_2457# a_n29_109# a_n287_n1197#
+ a_919_2545# a_1551_109# a_819_n1197# a_n129_n4851# a_819_4893# a_n1135_1327# a_n977_4981#
+ a_n1451_109# a_n1135_n3545# a_345_21# a_29_21# a_n1393_n1197# a_1293_n2415# a_603_n5981#
+ a_819_1239# a_n977_1327# a_n1609_n3545# a_n1077_4893# a_n1235_n4851# a_603_n2327#
+ a_n503_n3545# a_n29_3763# a_445_2545# a_n1077_1239# a_n503_109# a_n761_n1197# a_1235_n5981#
+ a_345_4893# a_187_n1197# a_1393_3763# a_n603_n4851# a_603_109# a_345_1239# a_1235_n2327#
+ a_1451_n1197# a_977_n2415# a_n761_2457# a_1293_2457# a_n919_4893# a_n503_4981# a_445_n5981#
+ a_129_4981# a_n1077_n4851# a_n129_n6069# a_n1293_4981# a_n919_1239# a_919_n5981#
+ a_n503_1327# a_n603_21# a_445_n2327# a_n345_n3545# a_661_n1197# a_129_1327# a_1077_n5981#
+ a_n187_3763# a_n1293_1327# a_1393_109# a_n819_n3545# a_977_4893# a_919_n2327# a_503_n4851#
+ a_n1293_109# a_n1235_n6069# a_n445_n4851# a_n1551_2457# a_1077_2545# a_n445_4893#
+ a_29_n3633# a_n1451_n3545# a_1077_n2327# a_977_1239# a_1293_n1197# a_n919_n4851#
+ a_n445_1239# a_1135_n4851# a_n1551_n4851# a_n603_n6069# a_287_n5981# a_n345_109#
+ a_29_3675# a_1551_n5981# a_287_n2327# a_n187_n3545# a_445_109# a_n1235_4893# a_1551_n2327#
+ a_345_n4851# a_977_n1197# a_n1077_n6069# a_n287_n4851# a_n1235_21# a_603_2545# a_n129_3675#
+ a_n1235_1239# a_n1293_n3545# a_503_4893# a_n661_4981# a_819_n4851# a_287_4981# a_761_n5981#
+ a_1551_3763# a_n29_n5981# a_503_n6069# a_503_1239# a_n661_1327# a_n1393_n4851# a_n445_n6069#
+ a_287_1327# a_761_n2327# a_n661_n3545# a_n819_3763# a_187_3675# a_n29_n2327# a_1451_2457#
+ a_503_21# a_n919_n6069# a_1393_n5981# a_1135_n6069# a_n1551_n6069# a_n761_n4851#
+ a_n1451_4981# a_1393_n2327# a_187_n4851# a_n345_3763# a_n1451_1327# a_1451_n4851#
+ a_n187_109# a_n1609_3763# a_1235_2545# a_n603_4893# a_345_n6069# a_n287_n6069# a_1135_4893#
+ a_287_109# a_n1393_4893# a_819_n6069# a_n603_1239# a_129_n4763# a_1135_1239# a_761_2545#
+ a_n977_n3545# a_661_n4851# a_n287_3675# a_n1393_1239# a_n1393_n6069# a_661_4893#
+ a_919_4981# a_129_n1109# a_n1135_3763# a_n1135_n5981# a_661_1239# a_919_1327# a_n129_n3633#
+ a_1293_n4851# a_819_3675# a_n977_3763# a_n1609_n5981# a_n761_n6069# a_n1135_n2327#
+ a_1135_21# a_187_n6069# a_n503_n5981# a_603_n4763# a_n919_21# a_n1609_n2327# a_445_4981#
+ a_n1077_3675# a_n1235_n3633# a_1451_n6069# a_603_n1109# a_n503_n2327# a_n761_21#
+ a_n1753_n6203# a_n29_2545# a_445_1327# a_345_3675# a_n129_21# a_1235_n4763# a_977_n4851#
+ a_n603_n3633# a_n761_4893# a_1393_2545# a_n819_109# a_1293_4893# a_1235_n1109# a_661_n6069#
+ a_919_109# a_n761_1239# a_1293_1239# a_n919_3675# a_n345_n5981# a_n503_3763# a_445_n4763#
+ a_129_3763# a_n1077_n3633# a_1293_n6069# a_n1293_3763# a_n819_n5981# a_919_n4763#
+ a_445_n1109# a_n345_n2327# a_1077_4981# a_n1551_4893# a_n1451_n5981# a_1077_n4763#
+ a_977_3675# a_n187_2545# a_919_n1109# a_n819_n2327# a_503_n3633# a_n445_n3633# a_n661_109#
+ a_n445_3675# a_n1551_1239# a_1077_1327# a_n1393_21# a_29_n2415# a_n1451_n2327# a_1077_n1109#
+ a_761_109# a_n919_n3633# a_1135_n3633# a_n1551_n3633# a_977_n6069# a_819_21# a_n187_n5981#
+ a_287_n4763# a_661_21# a_29_2457# a_n187_n2327# a_1551_n4763# a_287_n1109# a_603_4981#
+ a_n1235_3675# a_n1293_n5981# a_345_n3633# a_1551_n1109# a_n287_n3633# a_603_1327#
+ a_n129_2457# a_n1293_n2327# a_503_3675# a_n661_3763# a_819_n3633# a_287_3763# a_n661_n5981#
+ a_761_n4763# a_1551_2545# a_n29_n4763# a_1451_4893# a_n1393_n3633# a_n661_n2327#
+ a_761_n1109# a_n819_2545# a_187_2457# a_1451_1239# a_n29_n1109# a_1393_n4763# a_n761_n3633#
+ a_29_n1197# a_n1451_3763# a_187_n3633# a_1393_n1109# a_1235_4981# a_1451_n3633#
+ a_n345_2545# a_n603_3675# a_n1609_2545# a_1235_1327# a_1293_21# a_1135_3675# a_761_4981#
+ a_n977_n5981# a_n1393_3675# a_129_n3545# a_761_1327# a_n977_n2327# a_661_n3633#
+ a_n287_2457# a_661_3675# a_919_3763# a_n287_21# a_n1135_2545# a_n1135_n4763# a_1293_n3633#
X0 a_919_4981# a_819_4893# a_761_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_287_2545# a_187_2457# a_129_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X2 a_n1293_n5981# a_n1393_n6069# a_n1451_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X3 a_n661_109# a_n761_21# a_n819_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X4 a_n29_n5981# a_n129_n6069# a_n187_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X5 a_n187_n4763# a_n287_n4851# a_n345_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X6 a_1551_n5981# a_1451_n6069# a_1393_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X7 a_129_n2327# a_29_n2415# a_n29_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X8 a_n187_4981# a_n287_4893# a_n345_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X9 a_761_4981# a_661_4893# a_603_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X10 a_n1293_2545# a_n1393_2457# a_n1451_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X11 a_1393_2545# a_1293_2457# a_1235_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X12 a_129_109# a_29_21# a_n29_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X13 a_445_n1109# a_345_n1197# a_287_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X14 a_287_3763# a_187_3675# a_129_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X15 a_n187_109# a_n287_21# a_n345_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X16 a_n187_n5981# a_n287_n6069# a_n345_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X17 a_129_n3545# a_29_n3633# a_n29_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X18 a_n1293_3763# a_n1393_3675# a_n1451_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X19 a_1393_3763# a_1293_3675# a_1235_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X20 a_n345_1327# a_n445_1239# a_n503_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X21 a_445_n2327# a_345_n2415# a_287_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X22 a_287_4981# a_187_4893# a_129_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X23 a_919_n1109# a_819_n1197# a_761_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X24 a_n819_109# a_n919_21# a_n977_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X25 a_129_n4763# a_29_n4851# a_n29_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X26 a_n1293_4981# a_n1393_4893# a_n1451_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X27 a_1393_4981# a_1293_4893# a_1235_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X28 a_129_1327# a_29_1239# a_n29_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X29 a_n345_109# a_n445_21# a_n503_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X30 a_n345_2545# a_n445_2457# a_n503_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X31 a_445_n3545# a_345_n3633# a_287_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X32 a_1077_n1109# a_977_n1197# a_919_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X33 a_445_1327# a_345_1239# a_287_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X34 a_n1451_n1109# a_n1551_n1197# a_n1609_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X35 a_919_n2327# a_819_n2415# a_761_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X36 a_129_n5981# a_29_n6069# a_n29_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X37 a_129_2545# a_29_2457# a_n29_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X38 a_1551_1327# a_1451_1239# a_1393_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X39 a_n345_3763# a_n445_3675# a_n503_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X40 a_n1451_1327# a_n1551_1239# a_n1609_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X41 a_n503_109# a_n603_21# a_n661_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X42 a_445_n4763# a_345_n4851# a_287_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X43 a_1077_n2327# a_977_n2415# a_919_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X44 a_445_2545# a_345_2457# a_287_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X45 a_919_n3545# a_819_n3633# a_761_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X46 a_n1451_n2327# a_n1551_n2415# a_n1609_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X47 a_n345_n1109# a_n445_n1197# a_n503_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X48 a_129_3763# a_29_3675# a_n29_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X49 a_1551_2545# a_1451_2457# a_1393_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X50 a_n345_4981# a_n445_4893# a_n503_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X51 a_n1451_2545# a_n1551_2457# a_n1609_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X52 a_n29_109# a_n129_21# a_n187_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X53 a_445_n5981# a_345_n6069# a_287_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X54 a_1077_n3545# a_977_n3633# a_919_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X55 a_445_3763# a_345_3675# a_287_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X56 a_n977_1327# a_n1077_1239# a_n1135_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X57 a_919_n4763# a_819_n4851# a_761_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X58 a_n1451_n3545# a_n1551_n3633# a_n1609_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X59 a_n345_n2327# a_n445_n2415# a_n503_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X60 a_129_4981# a_29_4893# a_n29_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X61 a_1551_3763# a_1451_3675# a_1393_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X62 a_1077_1327# a_977_1239# a_919_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X63 a_1393_109# a_1293_21# a_1235_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X64 a_n1451_3763# a_n1551_3675# a_n1609_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X65 a_n503_1327# a_n603_1239# a_n661_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X66 a_n819_n1109# a_n919_n1197# a_n977_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X67 a_1077_n4763# a_977_n4851# a_919_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X68 a_445_4981# a_345_4893# a_287_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X69 a_n977_2545# a_n1077_2457# a_n1135_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X70 a_919_n5981# a_819_n6069# a_761_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X71 a_n1451_n4763# a_n1551_n4851# a_n1609_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X72 a_1077_109# a_977_21# a_919_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X73 a_n977_n1109# a_n1077_n1197# a_n1135_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X74 a_n345_n3545# a_n445_n3633# a_n503_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X75 a_1551_4981# a_1451_4893# a_1393_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X76 a_1077_2545# a_977_2457# a_919_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X77 a_n1451_4981# a_n1551_4893# a_n1609_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X78 a_n503_2545# a_n603_2457# a_n661_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X79 a_n819_n2327# a_n919_n2415# a_n977_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X80 a_1235_n1109# a_1135_n1197# a_1077_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X81 a_1551_109# a_1451_21# a_1393_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X82 a_1077_n5981# a_977_n6069# a_919_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X83 a_n977_3763# a_n1077_3675# a_n1135_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X84 a_603_1327# a_503_1239# a_445_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X85 a_n1451_n5981# a_n1551_n6069# a_n1609_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X86 a_n29_1327# a_n129_1239# a_n187_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X87 a_n345_n4763# a_n445_n4851# a_n503_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X88 a_n977_n2327# a_n1077_n2415# a_n1135_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X89 a_1077_3763# a_977_3675# a_919_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X90 a_1393_n1109# a_1293_n1197# a_1235_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X91 a_n503_3763# a_n603_3675# a_n661_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X92 a_n819_n3545# a_n919_n3633# a_n977_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X93 a_1235_n2327# a_1135_n2415# a_1077_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X94 a_761_109# a_661_21# a_603_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X95 a_603_n1109# a_503_n1197# a_445_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X96 a_n977_4981# a_n1077_4893# a_n1135_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X97 a_603_2545# a_503_2457# a_445_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X98 a_n29_2545# a_n129_2457# a_n187_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X99 a_n345_n5981# a_n445_n6069# a_n503_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X100 a_n977_n3545# a_n1077_n3633# a_n1135_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X101 a_1077_4981# a_977_4893# a_919_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X102 a_1393_n2327# a_1293_n2415# a_1235_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X103 a_n503_4981# a_n603_4893# a_n661_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X104 a_n819_n4763# a_n919_n4851# a_n977_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X105 a_1235_n3545# a_1135_n3633# a_1077_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X106 a_761_n1109# a_661_n1197# a_603_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X107 a_287_109# a_187_21# a_129_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X108 a_603_n2327# a_503_n2415# a_445_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X109 a_603_3763# a_503_3675# a_445_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X110 a_n1135_1327# a_n1235_1239# a_n1293_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X111 a_1235_1327# a_1135_1239# a_1077_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X112 a_1235_109# a_1135_21# a_1077_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X113 a_n29_3763# a_n129_3675# a_n187_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X114 a_n977_n4763# a_n1077_n4851# a_n1135_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X115 a_1393_n3545# a_1293_n3633# a_1235_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X116 a_919_109# a_819_21# a_761_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X117 a_n819_n5981# a_n919_n6069# a_n977_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X118 a_1235_n4763# a_1135_n4851# a_1077_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X119 a_761_n2327# a_661_n2415# a_603_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X120 a_603_n3545# a_503_n3633# a_445_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X121 a_445_109# a_345_21# a_287_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X122 a_603_4981# a_503_4893# a_445_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X123 a_n1135_2545# a_n1235_2457# a_n1293_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X124 a_1235_2545# a_1135_2457# a_1077_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X125 a_n29_4981# a_n129_4893# a_n187_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X126 a_n977_n5981# a_n1077_n6069# a_n1135_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X127 a_1393_n4763# a_1293_n4851# a_1235_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X128 a_1235_n5981# a_1135_n6069# a_1077_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X129 a_761_n3545# a_661_n3633# a_603_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X130 a_603_n4763# a_503_n4851# a_445_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X131 a_n1135_3763# a_n1235_3675# a_n1293_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X132 a_1235_3763# a_1135_3675# a_1077_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X133 a_603_109# a_503_21# a_445_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X134 a_n503_n1109# a_n603_n1197# a_n661_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X135 a_1393_n5981# a_1293_n6069# a_1235_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X136 a_761_n4763# a_661_n4851# a_603_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X137 a_603_n5981# a_503_n6069# a_445_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X138 a_287_n1109# a_187_n1197# a_129_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X139 a_n1135_4981# a_n1235_4893# a_n1293_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X140 a_1235_4981# a_1135_4893# a_1077_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X141 a_n503_n2327# a_n603_n2415# a_n661_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X142 a_n661_n1109# a_n761_n1197# a_n819_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X143 a_761_n5981# a_661_n6069# a_603_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X144 a_287_n2327# a_187_n2415# a_129_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X145 a_n1293_109# a_n1393_21# a_n1451_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X146 a_n1135_n1109# a_n1235_n1197# a_n1293_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X147 a_n503_n3545# a_n603_n3633# a_n661_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X148 a_n661_n2327# a_n761_n2415# a_n819_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X149 a_n819_1327# a_n919_1239# a_n977_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X150 a_287_n3545# a_187_n3633# a_129_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X151 a_n1293_n1109# a_n1393_n1197# a_n1451_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X152 a_n661_1327# a_n761_1239# a_n819_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X153 a_n503_n4763# a_n603_n4851# a_n661_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X154 a_n661_n3545# a_n761_n3633# a_n819_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X155 a_n1135_n2327# a_n1235_n2415# a_n1293_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X156 a_n29_n1109# a_n129_n1197# a_n187_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X157 a_n819_2545# a_n919_2457# a_n977_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X158 a_n1451_109# a_n1551_21# a_n1609_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X159 a_1551_n1109# a_1451_n1197# a_1393_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X160 a_287_n4763# a_187_n4851# a_129_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X161 a_919_1327# a_819_1239# a_761_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X162 a_n1293_n2327# a_n1393_n2415# a_n1451_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X163 a_n661_2545# a_n761_2457# a_n819_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X164 a_n503_n5981# a_n603_n6069# a_n661_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X165 a_n661_n4763# a_n761_n4851# a_n819_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X166 a_n1135_n3545# a_n1235_n3633# a_n1293_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X167 a_n29_n2327# a_n129_n2415# a_n187_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X168 a_n187_n1109# a_n287_n1197# a_n345_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X169 a_n819_3763# a_n919_3675# a_n977_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X170 a_n977_109# a_n1077_21# a_n1135_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X171 a_1551_n2327# a_1451_n2415# a_1393_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X172 a_n187_1327# a_n287_1239# a_n345_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X173 a_761_1327# a_661_1239# a_603_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X174 a_287_n5981# a_187_n6069# a_129_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X175 a_919_2545# a_819_2457# a_761_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X176 a_n1293_n3545# a_n1393_n3633# a_n1451_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X177 a_n661_3763# a_n761_3675# a_n819_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X178 a_n661_n5981# a_n761_n6069# a_n819_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X179 a_n1135_n4763# a_n1235_n4851# a_n1293_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X180 a_n29_n3545# a_n129_n3633# a_n187_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X181 a_n187_n2327# a_n287_n2415# a_n345_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X182 a_n819_4981# a_n919_4893# a_n977_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X183 a_1551_n3545# a_1451_n3633# a_1393_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X184 a_n187_2545# a_n287_2457# a_n345_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X185 a_761_2545# a_661_2457# a_603_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X186 a_n1135_109# a_n1235_21# a_n1293_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X187 a_919_3763# a_819_3675# a_761_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X188 a_n1293_n4763# a_n1393_n4851# a_n1451_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X189 a_n661_4981# a_n761_4893# a_n819_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X190 a_287_1327# a_187_1239# a_129_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X191 a_n1135_n5981# a_n1235_n6069# a_n1293_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X192 a_n29_n4763# a_n129_n4851# a_n187_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X193 a_n187_n3545# a_n287_n3633# a_n345_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X194 a_1551_n4763# a_1451_n4851# a_1393_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X195 a_129_n1109# a_29_n1197# a_n29_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X196 a_n187_3763# a_n287_3675# a_n345_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X197 a_761_3763# a_661_3675# a_603_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X198 a_n1293_1327# a_n1393_1239# a_n1451_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X199 a_1393_1327# a_1293_1239# a_1235_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6 a_n108_n250# w_n308_n547# a_50_n250# a_n50_n347#
X0 a_50_n250# a_n50_n347# a_n108_n250# w_n308_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0 a_50_n200# a_n108_n200# a_n50_n288# a_n252_n422#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n252_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_L9TFKV a_n958_n300# a_n900_n388# a_n1092_n522#
+ a_900_n300#
X0 a_900_n300# a_n900_n388# a_n958_n300# a_n1092_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=9
.ends

.subckt sky130_am_ip__ldo_01v8 AVDD VOUT AVSS ENA VREF_EXT SEL_EXT DVDD DVSS
XXM56 vbias_p vy AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM67 vbias_n vbias_n vbias_n vbias_n AVSS AVSS vbias_n AVSS vbias_n vbias_n vbias_n
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM78 AVSS AVSS nena ena_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM89 AVSS verr AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM46 vbias_p vx AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM57 vbias_c verr AVDD vy sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM68 AVDD vbias_c vbias_c AVDD sky130_fd_pr__pfet_g5v0d10v5_PC2PN5
XXM79 vbias_p vref_int AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
Xx1 ENA DVDD DVSS AVDD AVDD ena_3v3 AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
XXM58 vbias_c m2_8539_n7649# AVDD vx sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM69 vbias_n vbias_n vbias_c vbias_n AVSS AVSS vbias_c AVSS vbias_c vbias_c vbias_c
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
Xx2 SEL_EXT DVDD DVSS AVDD AVDD sel_ext_3v3 AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
XXM48 verr AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXM59 verr AVSS AVDD vpass sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXR4 m1_5119_3142# m1_5119_2478# m1_5119_1150# m1_7519_2644# m1_7519_984# m1_7519_1980#
+ m1_5119_2146# m1_5119_3474# m1_7519_1648# m1_5119_1482# m1_7519_2976# m1_5119_2810#
+ vm m1_7519_2976# m1_5119_818# m1_5119_1814# m1_5119_1482# m1_7519_1316# m1_5119_3474#
+ m1_7519_3308# m1_5119_3142# m1_5119_2146# m1_7519_1648# m1_7519_2312# m1_7519_2644#
+ VOUT m1_5119_1150# AVSS m1_5119_2478# m1_7519_1316# m1_5119_2810# m1_7519_3308#
+ m1_7519_2312# m1_5119_818# m1_7519_1980# m1_5119_1814# m1_7519_984# sky130_fd_pr__res_xhigh_po_0p35_QZEXQH
XXR5 m1_5117_n1479# m1_5117_n2475# m1_7517_n4965# m1_5117_n4799# m1_7517_n981# m1_5117_n3803#
+ m1_5117_181# m1_7517_n1977# m1_7517_n3637# m1_7517_n2641# m1_7517_n4633# m1_5117_n815#
+ m1_7517_15# m1_5117_n2475# m1_5117_n5463# m1_5117_n151# m1_5117_n4467# m1_7517_n649#
+ m1_5117_n3471# m1_7517_n2973# m1_5117_n1147# vm m1_7517_n1645# m1_5117_181# m1_5117_n2143#
+ m1_7517_n3969# m1_7517_n4965# m1_5117_n815# m1_5117_n5131# m1_5117_n4135# m1_7517_n1977#
+ m1_5117_n2807# m1_7517_n981# m1_5117_n483# m1_7517_15# m1_7517_n3305# m1_5117_n3139#
+ m1_7517_n4301# m1_7517_n5297# m1_5117_n1479# m1_7517_n1645# m1_7517_n649# m1_7517_n4301#
+ m1_5117_n1811# m1_5117_n2807# m1_7517_n3305# m1_5117_n5463# m1_7517_n5297# m1_5117_n4467#
+ m1_7517_n2641# m1_5117_n151# m1_7517_n2309# m1_7517_n1313# m1_5117_n3471# m1_7517_n317#
+ m1_7517_n4633# m1_5117_n2143# m1_5117_n4799# m1_7517_n3637# AVSS AVSS m1_5117_n1147#
+ m1_5117_n1811# m1_5117_n5131# m1_7517_n1313# m1_5117_n3803# m1_7517_n2309# m1_5117_n483#
+ m1_5117_n4135# m1_7517_n3969# m1_7517_n317# m1_5117_n3139# m1_7517_n2973# sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H
XXR6 AVSS m1_22164_n7435# AVSS m1_22164_n7435# m2_26640_n7437# sky130_fd_pr__res_xhigh_po_0p35_743D3R
XXC1[0] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[1] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[2] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC3 AVSS vref sky130_fd_pr__cap_mim_m3_1_VCAG9S__0
XXM90 nena vdd_start AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM80 vref_int AVSS m1_12626_n9400# m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM70 AVSS vdd_start vbias_n vstart sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM81 vref_int AVSS vref_int m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM60 vbias_p vpass AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM71 m1_20910_n7332# vstart vstart AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM82 vref_int AVSS m1_12626_n9400# AVSS sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM72 m1_20184_n7334# m1_20910_n7332# m1_20910_n7332# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM83 AVSS AVSS nsel_ext sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM61[0] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[1] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[2] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[3] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[4] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM62 vbias_p AVDD AVDD m1_19028_n7338# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM73 AVDD m1_20184_n7334# m1_20184_n7334# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM84 AVDD AVDD nsel_ext sel_ext_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
Xsky130_fd_pr__pfet_g5v0d10v5_KLAZY6_0 ena_3v3 vbias_c AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM52 vy m2_6784_n8214# vm AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM63 vbias_c m1_19028_n7338# AVDD vbias_p sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM74 vbias_n vbias_n vstart vbias_n AVSS AVSS vstart AVSS vstart vstart vstart vbias_n
+ AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM85 AVSS vbias_n AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM53 vx m2_6784_n8214# vref AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM64 vbias_p AVDD AVDD m1_16878_n7330# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM75 AVSS vref vref_int nsel_ext sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM54 AVSS vbias_n AVSS m2_6784_n8214# sky130_fd_pr__nfet_g5v0d10v5_L9TFKV
XXM65 vbias_c m1_16878_n7330# AVDD vbias_n sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM76 AVDD AVDD nena ena_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
XXM87 AVSS vpass AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM55 m2_8539_n7649# AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXM66[0] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[1] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[2] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[3] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM77 AVSS VREF_EXT vref sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM88 ena_3v3 vbias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_QTPFY2 a_n29_n1250# a_n945_n1250# a_n429_n1338# a_945_n1338#
+ a_n487_n1250# a_n887_n1338# a_1803_n1250# a_487_n1338# a_1345_n1250# a_n1963_n1424#
+ a_n1403_n1250# a_n1803_n1338# a_429_n1250# a_n1861_n1250# a_887_n1250# a_n1345_n1338#
+ a_1403_n1338# a_29_n1338#
X0 a_n487_n1250# a_n887_n1338# a_n945_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X1 a_n945_n1250# a_n1345_n1338# a_n1403_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X2 a_887_n1250# a_487_n1338# a_429_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X3 a_1803_n1250# a_1403_n1338# a_1345_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=2
X4 a_1345_n1250# a_945_n1338# a_887_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X5 a_n1403_n1250# a_n1803_n1338# a_n1861_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=2
X6 a_n29_n1250# a_n429_n1338# a_n487_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X7 a_429_n1250# a_29_n1338# a_n29_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_QGRVRG a_n360_n674# a_200_n500# a_n258_n500# a_n200_n588#
X0 a_200_n500# a_n200_n588# a_n258_n500# a_n360_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__nfet_01v8_ME6MQD a_1000_n1000# a_n1160_n1174# a_n1000_n1088#
+ a_n1058_n1000#
X0 a_1000_n1000# a_n1000_n1088# a_n1058_n1000# a_n1160_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_6H4ZLK a_n1000_n597# a_1000_n500# a_n1058_n500# w_n1196_n719#
X0 a_1000_n500# a_n1000_n597# a_n1058_n500# w_n1196_n719# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_D2R37Y a_1000_n500# a_n1058_n500# a_n1000_n588# a_n1160_n674#
X0 a_1000_n500# a_n1000_n588# a_n1058_n500# a_n1160_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_5TKQ2R a_500_n1000# a_n660_n1174# a_n500_n1088# a_n558_n1000#
X0 a_500_n1000# a_n500_n1088# a_n558_n1000# a_n660_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=5
.ends

.subckt sbvfcm vdd pbias nbias vx vss XM7/w_n1196_n719# XM8/w_n1196_n719# VSUBS
Xsky130_fd_pr__nfet_01v8_QTPFY2_0 m1_5880_1010# m1_5880_1010# m1_5868_n3400# m1_5868_n3400#
+ vx m1_5868_n3400# m1_5880_1010# m1_5868_n3400# vx VSUBS vx m1_5868_n3400# vx m1_5880_1010#
+ m1_5880_1010# m1_5868_n3400# m1_5868_n3400# m1_5868_n3400# sky130_fd_pr__nfet_01v8_QTPFY2
XXM4 VSUBS m1_9368_n812# vss m1_5868_n3400# sky130_fd_pr__nfet_01v8_QGRVRG
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0 m1_9568_n2160# vdd sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM5 pbias VSUBS nbias m1_5880_1010# sky130_fd_pr__nfet_01v8_ME6MQD
XXM6 m1_9368_n812# VSUBS nbias m1_5868_n3400# sky130_fd_pr__nfet_01v8_ME6MQD
XXM7 pbias pbias vdd XM7/w_n1196_n719# sky130_fd_pr__pfet_01v8_6H4ZLK
XXM8 pbias vdd m1_5868_n3400# XM8/w_n1196_n719# sky130_fd_pr__pfet_01v8_6H4ZLK
XXC1 m1_9568_n2160# vdd sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM10 pbias vss m1_9568_n2160# VSUBS sky130_fd_pr__nfet_01v8_D2R37Y
XXM11 vss VSUBS m1_5868_n3400# m1_9568_n2160# sky130_fd_pr__nfet_01v8_5TKQ2R
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_H5FMR6 a_n199_n891# a_n69_n761# a_n69_329#
X0 a_n69_329# a_n69_n761# a_n199_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_H5TM75 a_n420_n761# a_n550_n891# a_n420_329#
+ a_48_n761# a_n186_n761# a_282_329# a_48_329# a_n186_329# a_282_n761#
X0 a_n420_329# a_n420_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_48_329# a_48_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X2 a_282_329# a_282_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X3 a_n186_329# a_n186_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__nfet_01v8_J222PV a_n429_n588# a_29_n588# a_n589_n674# a_n487_n500#
+ a_n29_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_D5BT6X a_n420_n761# a_n654_329# a_n888_329#
+ a_n420_329# a_48_n761# a_n654_n761# a_n1018_n891# a_n888_n761# a_n186_n761# a_750_n761#
+ a_282_329# a_48_329# a_n186_329# a_282_n761# a_750_329# a_516_n761# a_516_329#
X0 a_n420_329# a_n420_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_48_329# a_48_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X2 a_282_329# a_282_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X3 a_n888_329# a_n888_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X4 a_750_329# a_750_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X5 a_516_329# a_516_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X6 a_n186_329# a_n186_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X7 a_n654_329# a_n654_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_2G52HS a_48_n761# a_n186_n761# a_n316_n891#
+ a_48_329# a_n186_329#
X0 a_48_329# a_48_n761# a_n316_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_n186_329# a_n186_n761# a_n316_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt trim_res A trim0 trim2 trim3 trim1 B VSUBS
Xsky130_fd_pr__res_xhigh_po_0p69_H5FMR6_0 VSUBS m1_835_n1590# B sky130_fd_pr__res_xhigh_po_0p69_H5FMR6
Xsky130_fd_pr__res_xhigh_po_0p69_H5TM75_0 m1_834_n3490# VSUBS m1_4520_n760# m1_4760_n1840#
+ m1_4760_n1840# m1_4980_n760# m1_4980_n760# m1_4520_n760# m1_1200_n3120# sky130_fd_pr__res_xhigh_po_0p69_H5TM75
XXM1 trim0 trim0 VSUBS B m1_835_n1590# B sky130_fd_pr__nfet_01v8_J222PV
XXM2 trim1 trim1 VSUBS m1_835_n1590# m1_834_n3490# m1_835_n1590# sky130_fd_pr__nfet_01v8_J222PV
XXM3 trim2 trim2 VSUBS m1_834_n3490# m1_1200_n3120# m1_834_n3490# sky130_fd_pr__nfet_01v8_J222PV
XXM4 trim3 trim3 VSUBS m1_1200_n3120# A m1_1200_n3120# sky130_fd_pr__nfet_01v8_J222PV
Xsky130_fd_pr__res_xhigh_po_0p69_D5BT6X_0 m1_4020_n3720# m1_3780_n2640# A m1_3780_n2640#
+ m1_4500_n3720# m1_3560_n3720# VSUBS m1_3560_n3720# m1_4020_n3720# m1_4960_n3720#
+ m1_4720_n2640# m1_4260_n2640# m1_4260_n2640# m1_4500_n3720# m1_1200_n3120# m1_4960_n3720#
+ m1_4720_n2640# sky130_fd_pr__res_xhigh_po_0p69_D5BT6X
Xsky130_fd_pr__res_xhigh_po_0p69_2G52HS_0 m1_834_n3490# m1_835_n1590# VSUBS m1_3920_n760#
+ m1_3920_n760# sky130_fd_pr__res_xhigh_po_0p69_2G52HS
.ends

.subckt sky130_fd_pr__nfet_01v8_QGMQL3 a_n158_n250# a_n100_n338# a_n260_n424# a_100_n250#
X0 a_100_n250# a_n100_n338# a_n158_n250# a_n260_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_MMMA4V a_100_n500# a_n158_n500# a_n100_n588# a_n260_n674#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_HS3BL4 a_100_n800# a_n158_n800# a_n100_n888# a_n260_n974#
X0 a_100_n800# a_n100_n888# a_n158_n800# a_n260_n974# sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_W2FWA4 a_n429_n588# a_29_n588# a_n589_n674# a_n487_n500#
+ a_n29_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_ST5LSM a_n1087_n2000# w_n1225_n2219# a_n1029_n2097#
+ a_n29_n2000# a_1029_n2000# a_29_n2097#
X0 a_n29_n2000# a_n1029_n2097# a_n1087_n2000# w_n1225_n2219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
X1 a_1029_n2000# a_29_n2097# a_n29_n2000# w_n1225_n2219# sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_CXW7PW a_n487_n1000# a_429_n1000# a_29_n1088#
+ a_n621_n1222# a_n429_n1088# a_n29_n1000#
X0 a_429_n1000# a_29_n1088# a_n29_n1000# a_n621_n1222# sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=2
X1 a_n29_n1000# a_n429_n1088# a_n487_n1000# a_n621_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=2
.ends

.subckt output_amp vo vp vn ibias vss vdd VSUBS
XXM1 ibias ibias VSUBS vss sky130_fd_pr__nfet_01v8_QGMQL3
XXM2 vss vcm ibias VSUBS sky130_fd_pr__nfet_01v8_MMMA4V
XXM3 vo vss ibias VSUBS sky130_fd_pr__nfet_01v8_HS3BL4
XXM4 vn vn VSUBS vcm m1_5267_n942# vcm sky130_fd_pr__nfet_01v8_W2FWA4
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[0] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[1] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[2] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[3] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[4] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM5 vp vp VSUBS vcm m1_7167_n942# vcm sky130_fd_pr__nfet_01v8_J222PV
XXM6 m1_5168_2580# vdd m1_5168_2580# vdd sky130_fd_pr__pfet_01v8_6H4ZLK
XXM7 m1_5168_2580# vo_pre vdd vdd sky130_fd_pr__pfet_01v8_6H4ZLK
XXM8 vdd vdd vo_pre vo vdd vo_pre sky130_fd_pr__pfet_01v8_ST5LSM
XXM9 m1_5267_n942# m1_5267_n942# vn VSUBS vn m1_5168_2580# sky130_fd_pr__nfet_05v0_nvt_CXW7PW
XXC2[0] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[1] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[2] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[3] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[4] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM10 m1_7167_n942# m1_7167_n942# vp VSUBS vp vo_pre sky130_fd_pr__nfet_05v0_nvt_CXW7PW
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_E9MCU4 a_n433_n2363# a_n69_n2233# a_n69_1801#
+ a_165_1801# a_165_n2233# a_n303_n2233# a_n303_1801#
X0 a_n69_1801# a_n69_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
X1 a_165_1801# a_165_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
X2 a_n303_1801# a_n303_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_39QBTQ a_n69_844# a_n69_n1276# a_n199_n1406#
X0 a_n69_844# a_n69_n1276# a_n199_n1406# sky130_fd_pr__res_xhigh_po_0p69 l=8.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH a_n420_1847# a_n186_n2279# a_n550_n2409#
+ a_48_1847# a_n186_1847# a_282_n2279# a_48_n2279# a_n420_n2279# a_282_1847#
X0 a_n186_1847# a_n186_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X1 a_n420_1847# a_n420_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X2 a_48_1847# a_48_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X3 a_282_1847# a_282_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_GAZAU4 a_984_n2306# a_n186_1874# a_750_1874#
+ a_n1590_1874# a_984_1874# a_n1590_n2306# a_1218_n2306# a_282_n2306# a_n1720_n2436#
+ a_282_1874# a_48_n2306# a_n420_n2306# a_n1122_1874# a_1218_1874# a_750_n2306# a_516_1874#
+ a_n1356_1874# a_n1356_n2306# a_n420_1874# a_n888_n2306# a_516_n2306# a_48_1874#
+ a_n654_1874# a_n1122_n2306# a_n186_n2306# a_n888_1874# a_1452_n2306# a_1452_1874#
+ a_n654_n2306#
X0 a_n654_1874# a_n654_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X1 a_n186_1874# a_n186_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X2 a_516_1874# a_516_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X3 a_n420_1874# a_n420_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X4 a_1452_1874# a_1452_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X5 a_n1590_1874# a_n1590_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X6 a_48_1874# a_48_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X7 a_984_1874# a_984_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X8 a_n1356_1874# a_n1356_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X9 a_1218_1874# a_1218_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X10 a_750_1874# a_750_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X11 a_n1122_1874# a_n1122_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X12 a_n888_1874# a_n888_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X13 a_282_1874# a_282_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
.ends

.subckt sky130_fd_pr__nfet_01v8_2333C8 a_n2000_n338# a_n2160_n424# a_2000_n250# a_n2058_n250#
X0 a_2000_n250# a_n2000_n338# a_n2058_n250# a_n2160_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_Q33MQV a_1000_n200# a_n1058_n200# a_n1000_n288# a_n1160_n374#
X0 a_1000_n200# a_n1000_n288# a_n1058_n200# a_n1160_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=10
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_B3G3L7 a_n29_n2618# a_n2029_21# a_29_21# w_n2225_n2837#
+ a_2029_118# a_2029_n2618# a_n2029_n2715# a_29_n2715# a_n2087_118# a_n29_118# a_n2087_n2618#
X0 a_2029_118# a_29_21# a_n29_118# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=10
X1 a_n29_118# a_n2029_21# a_n2087_118# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=10
X2 a_n29_n2618# a_n2029_n2715# a_n2087_n2618# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=10
X3 a_2029_n2618# a_29_n2715# a_n29_n2618# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=10
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_pr__pfet_01v8_XPMKX6 a_30_n1000# a_n33_n1097# a_n88_n1000# w_n226_n1219#
X0 a_30_n1000# a_n33_n1097# a_n88_n1000# w_n226_n1219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.3
.ends

.subckt sky130_ak_ip__cmos_vref vbg avdd18 ena vbgsc vbgtg trim3 trim2 trim1 trim0
+ vptat dvdd avss dvss
Xsky130_fd_sc_hd__buf_1_4 trim1 dvss dvss dvdd dvdd trim1buf sky130_fd_sc_hd__buf_1
Xx1 avdd_ena pbias vref vptat avss avdd_ena avdd_ena avss sbvfcm
Xx3 x3/A trim0buf trim2buf trim3buf trim1buf avss avss trim_res
Xx2 vbg vref x2/vn x2/ibias avss avdd_ena avss output_amp
XR1 avss m1_9471_n10626# m1_9471_n10158# vbgtg m1_9471_n10626# m1_9471_n10158# vbg
+ sky130_fd_pr__res_xhigh_po_0p69_E9MCU4
XR2 vbgtg vbgsc avss sky130_fd_pr__res_xhigh_po_0p69_39QBTQ
XR3 vbgsc m1_9472_n11356# avss m1_13592_n11600# m1_13592_n11600# m1_9472_n11824# m1_9472_n11824#
+ m1_9472_n11356# x2/vn sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH
XR4 m1_13651_n12750# m1_9472_n13920# m1_9472_n12984# m1_9472_n15324# m1_9472_n12984#
+ x3/A m1_13651_n12750# m1_13651_n13686# avss m1_9472_n13452# m1_13651_n13686# m1_13651_n14154#
+ m1_9472_n14856# m1_9472_n12516# m1_13651_n13218# m1_9472_n13452# m1_9472_n15324#
+ m1_13651_n15090# m1_9472_n14388# m1_13651_n14622# m1_13651_n13218# m1_9472_n13920#
+ m1_9472_n14388# m1_13651_n15090# m1_13651_n14154# m1_9472_n14856# x2/vn m1_9472_n12516#
+ m1_13651_n14622# sky130_fd_pr__res_xhigh_po_0p69_GAZAU4
XXM1 vref avss vptat avss sky130_fd_pr__nfet_01v8_2333C8
XXM2 vptat vref vref avss sky130_fd_pr__nfet_01v8_Q33MQV
Xsky130_fd_sc_hd__inv_2_0 ena dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2
XXM3 pbias x2/ibias avdd_ena avdd_ena sky130_fd_pr__pfet_01v8_6H4ZLK
Xsky130_fd_sc_hd__diode_2_0 trim2 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
XXM9 vref pbias pbias avdd_ena avdd_ena avdd_ena pbias pbias avdd_ena vref avdd_ena
+ sky130_fd_pr__pfet_01v8_B3G3L7
Xsky130_fd_sc_hd__diode_2_1 ena dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_2 trim3 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_3 trim1 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_6_0 dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__diode_2_4 trim0 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_1_0 trim0 dvss dvss dvdd dvdd trim0buf sky130_fd_sc_hd__buf_1
XXM20 avdd_ena sky130_fd_sc_hd__inv_2_0/Y avdd18 dvdd sky130_fd_pr__pfet_01v8_XPMKX6
Xsky130_fd_sc_hd__buf_1_2 trim3 dvss dvss dvdd dvdd trim3buf sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 trim2 dvss dvss dvdd dvdd trim2buf sky130_fd_sc_hd__buf_1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7 a_n445_n1088# a_n503_n1000# a_345_n1088#
+ a_n287_n1088# a_n345_n1000# a_187_n1088# a_n187_n1000# a_129_n1000# a_29_n1088#
+ a_445_n1000# a_287_n1000# a_n129_n1088# a_n637_n1222# a_n29_n1000#
X0 a_445_n1000# a_345_n1088# a_287_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n29_n1000# a_n129_n1088# a_n187_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n187_n1000# a_n287_n1088# a_n345_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_287_n1000# a_187_n1088# a_129_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n345_n1000# a_n445_n1088# a_n503_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 a_129_n1000# a_29_n1088# a_n29_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQSWZU a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_29_n1097# a_n187_n1000# a_n661_n1000# a_n977_n1000# a_n129_n1097# a_n603_n1097#
+ a_503_n1097# a_n445_n1097# a_n919_n1097# a_345_n1097# a_n287_n1097# a_819_n1097#
+ a_187_n1097# a_n761_n1097# w_n1177_n1297# a_129_n1000# a_661_n1097# a_603_n1000#
+ a_919_n1000# a_445_n1000# a_287_n1000# a_761_n1000# a_n29_n1000#
X0 a_129_n1000# a_29_n1097# a_n29_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_445_n1000# a_345_n1097# a_287_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n503_n1000# a_n603_n1097# a_n661_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n29_n1000# a_n129_n1097# a_n187_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_603_n1000# a_503_n1097# a_445_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 a_n819_n1000# a_n919_n1097# a_n977_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X6 a_n661_n1000# a_n761_n1097# a_n819_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 a_919_n1000# a_819_n1097# a_761_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X8 a_n187_n1000# a_n287_n1097# a_n345_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_761_n1000# a_661_n1097# a_603_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X10 a_287_n1000# a_187_n1097# a_129_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X11 a_n345_n1000# a_n445_n1097# a_n503_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt isolated_switch_4 on off in vdd shunt out vss
XXM15 on m2_961_n2337# on on out on m2_961_n2337# m2_961_n2337# on m2_961_n2337# out
+ on vss out sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7
XXM4 m2_961_n2337# out m2_961_n2337# off m2_961_n2337# out out off off off off off
+ off off off off off vdd m2_961_n2337# off out out m2_961_n2337# out m2_961_n2337#
+ out sky130_fd_pr__pfet_g5v0d10v5_AQSWZU
Xsky130_fd_pr__nfet_g5v0d10v5_F5JQJ7_0 on in on on m2_961_n2337# on in in on in m2_961_n2337#
+ on vss m2_961_n2337# sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7
Xsky130_fd_pr__nfet_g5v0d10v5_EJGQJV_0 vss vss m2_961_n2337# shunt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
Xsky130_fd_pr__pfet_g5v0d10v5_AQSWZU_0 in m2_961_n2337# in off in m2_961_n2337# m2_961_n2337#
+ off off off off off off off off off off vdd in off m2_961_n2337# m2_961_n2337# in
+ m2_961_n2337# in m2_961_n2337# sky130_fd_pr__pfet_g5v0d10v5_AQSWZU
.ends

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
.ends

.subckt isolated_switch_xlarge on out in avdd off avss dvdd dvss
Xx2 on dvdd dvss avdd avdd x2/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xx3 off dvdd dvss avdd avdd x3/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xisolated_switch_4_0 x2/X isolated_switch_4_0/off in avdd x3/X out avss isolated_switch_4
Xsky130_fd_sc_hvl__diode_2_0 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_1 off dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_1_0 x2/X dvss dvss avdd avdd isolated_switch_4_0/off sky130_fd_sc_hvl__inv_1
.ends

.subckt switch_array_2 channel0_in_to_out[1] channel0_in_to_out[0] channel1_in_to_out[1]
+ channel1_in_to_out[0] channel0_in channel0_out channel1_in channel1_out avdd dvdd
+ avss dvss
Xisolated_switch_xlarge_0[0] channel1_in_to_out[0] channel1_out channel1_in avdd channel1_in_to_out[1]
+ avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[1] channel0_in_to_out[0] channel0_out channel0_in avdd channel0_in_to_out[1]
+ avss dvdd dvss isolated_switch_xlarge
.ends

.subckt ct2_switch_array switch_array_2_0/dvdd switch_array_2_0/channel0_in switch_array_2_0/channel1_in_to_out[1]
+ switch_array_2_0/channel1_in_to_out[0] switch_array_2_0/channel1_out switch_array_2_0/avdd
+ switch_array_2_0/avss switch_array_2_0/channel0_in_to_out[1] switch_array_2_0/channel0_in_to_out[0]
+ switch_array_2_0/channel1_in VSUBS
Xswitch_array_2_0 switch_array_2_0/channel0_in_to_out[1] switch_array_2_0/channel0_in_to_out[0]
+ switch_array_2_0/channel1_in_to_out[1] switch_array_2_0/channel1_in_to_out[0] switch_array_2_0/channel0_in
+ switch_array_2_0/channel1_out switch_array_2_0/channel1_in switch_array_2_0/channel1_out
+ switch_array_2_0/avdd switch_array_2_0/dvdd switch_array_2_0/avss VSUBS switch_array_2
.ends

.subckt audiodac_drv_latch in_p in_n vdd_hi vss
X0 in_p in_n vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X1 vss in_p in_n vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X2 in_n in_p vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X3 vdd_hi in_n in_p vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X4 in_p in_n vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 vdd_hi in_p in_n vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X6 in_n in_p vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X7 vss in_n in_p vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CYU746 a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_29_n1097# a_n187_n1000# a_n661_n1000# a_n129_n1097# a_n603_n1097# w_n1019_n1297#
+ a_503_n1097# a_n445_n1097# a_345_n1097# a_n287_n1097# a_187_n1097# a_n761_n1097#
+ a_129_n1000# a_661_n1097# a_603_n1000# a_445_n1000# a_287_n1000# a_761_n1000# a_n29_n1000#
X0 a_129_n1000# a_29_n1097# a_n29_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_445_n1000# a_345_n1097# a_287_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n503_n1000# a_n603_n1097# a_n661_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n29_n1000# a_n129_n1097# a_n187_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_603_n1000# a_503_n1097# a_445_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 a_n661_n1000# a_n761_n1097# a_n819_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X6 a_n187_n1000# a_n287_n1097# a_n345_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 a_761_n1000# a_661_n1097# a_603_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X8 a_287_n1000# a_187_n1097# a_129_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_n345_n1000# a_n445_n1097# a_n503_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QABAEG a_30_n588# a_288_n500# a_n478_n722# a_n128_n588#
+ a_188_n588# a_n286_n588# a_130_n500# a_n28_n500# a_n186_n500# a_n344_n500#
X0 a_n28_n500# a_n128_n588# a_n186_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_288_n500# a_188_n588# a_130_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X2 a_n186_n500# a_n286_n588# a_n344_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X3 a_130_n500# a_30_n588# a_n28_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3 a_n242_n622# a_50_n400# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n242_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YSH3F7 a_503_n1088# a_n445_n1088# a_n953_n1222#
+ a_n503_n1000# a_345_n1088# a_n287_n1088# a_n345_n1000# a_n819_n1000# a_187_n1088#
+ a_n761_n1088# a_n187_n1000# a_661_n1088# a_n661_n1000# a_129_n1000# a_29_n1088#
+ a_603_n1000# a_445_n1000# a_287_n1000# a_n129_n1088# a_761_n1000# a_n29_n1000# a_n603_n1088#
X0 a_445_n1000# a_345_n1088# a_287_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n503_n1000# a_n603_n1088# a_n661_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n29_n1000# a_n129_n1088# a_n187_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_603_n1000# a_503_n1088# a_445_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n661_n1000# a_n761_n1088# a_n819_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 a_n187_n1000# a_n287_n1088# a_n345_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 a_761_n1000# a_661_n1088# a_603_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X7 a_287_n1000# a_187_n1088# a_129_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X8 a_n345_n1000# a_n445_n1088# a_n503_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_129_n1000# a_29_n1088# a_n29_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QCNVDG a_n108_n1000# a_n366_n1088# a_n424_n1000#
+ a_266_n1088# a_n266_n1000# a_50_n1000# a_208_n1000# a_366_n1000# a_n50_n1088# a_n208_n1088#
+ a_108_n1088# a_n558_n1222#
X0 a_n266_n1000# a_n366_n1088# a_n424_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X1 a_366_n1000# a_266_n1088# a_208_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X2 a_50_n1000# a_n50_n1088# a_n108_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n108_n1000# a_n208_n1088# a_n266_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_208_n1000# a_108_n1088# a_50_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WECJAU a_30_n1098# a_n28_n1000# a_n344_n1000#
+ a_n186_n1000# a_130_n1000# a_188_n1098# a_n128_n1098# a_288_n1000# a_n286_n1098#
+ w_n544_n1296#
X0 a_130_n1000# a_30_n1098# a_n28_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n28_n1000# a_n128_n1098# a_n186_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_288_n1000# a_188_n1098# a_130_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n186_n1000# a_n286_n1098# a_n344_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_54K6JW a_445_118# a_n345_118# a_n661_n2118# a_n187_118#
+ a_187_21# a_287_118# a_n445_21# a_n819_118# a_n661_118# a_761_118# a_345_21# a_29_21#
+ a_n603_21# a_129_n2118# a_29_n2215# a_603_n2118# a_503_21# a_445_n2118# a_287_n2118#
+ a_n129_n2215# a_761_n2118# a_n29_n2118# a_129_118# a_n129_21# a_n761_21# a_n603_n2215#
+ w_n1019_n2415# a_503_n2215# a_n445_n2215# a_n29_118# a_661_21# a_n503_n2118# a_345_n2215#
+ a_n287_n2215# a_603_118# a_n503_118# a_n345_n2118# a_187_n2215# a_n761_n2215# a_n819_n2118#
+ a_n187_n2118# a_661_n2215# a_n287_21#
X0 a_603_118# a_503_21# a_445_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_287_n2118# a_187_n2215# a_129_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n661_n2118# a_n761_n2215# a_n819_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X3 a_n29_n2118# a_n129_n2215# a_n187_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n187_n2118# a_n287_n2215# a_n345_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 a_129_n2118# a_29_n2215# a_n29_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 a_445_n2118# a_345_n2215# a_287_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 a_n661_118# a_n761_21# a_n819_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X8 a_129_118# a_29_21# a_n29_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_n187_118# a_n287_21# a_n345_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X10 a_n345_118# a_n445_21# a_n503_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X11 a_n503_118# a_n603_21# a_n661_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X12 a_n345_n2118# a_n445_n2215# a_n503_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X13 a_n29_118# a_n129_21# a_n187_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X14 a_603_n2118# a_503_n2215# a_445_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X15 a_761_118# a_661_21# a_603_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X16 a_761_n2118# a_661_n2215# a_603_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X17 a_287_118# a_187_21# a_129_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X18 a_445_118# a_345_21# a_287_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X19 a_n503_n2118# a_n603_n2215# a_n661_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HKUKAU a_30_n162# w_n386_n362# a_n28_n64# a_n128_n162#
+ a_n186_n64# a_130_n64#
X0 a_n28_n64# a_n128_n162# a_n186_n64# w_n386_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_130_n64# a_30_n162# a_n28_n64# w_n386_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3QQKN5 a_130_n400# w_n386_n696# a_n28_n400# a_n186_n400#
+ a_n128_n498# a_30_n498#
X0 a_n28_n400# a_n128_n498# a_n186_n400# w_n386_n696# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_130_n400# a_30_n498# a_n28_n400# w_n386_n696# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt audiodac_drv_lite_half in crosscon out vdd_hi vss
Xsky130_fd_pr__pfet_g5v0d10v5_CYU746_0 vdd_hi drv4 vdd_hi crosscon vdd_hi drv4 crosscon
+ crosscon vdd_hi crosscon crosscon crosscon crosscon crosscon crosscon vdd_hi crosscon
+ drv4 vdd_hi drv4 vdd_hi drv4 sky130_fd_pr__pfet_g5v0d10v5_CYU746
Xsky130_fd_pr__nfet_g5v0d10v5_QABAEG_0 drv2 vss vss drv2 drv2 drv2 crosscon vss crosscon
+ vss sky130_fd_pr__nfet_g5v0d10v5_QABAEG
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ3_0 vss drv2 vss drv1 sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
Xsky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0 vss vss drv1 in sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ
Xsky130_fd_pr__nfet_g5v0d10v5_YSH3F7_0 drv4 drv4 vss vss drv4 drv4 out vss drv4 drv4
+ vss drv4 out vss drv4 out vss out drv4 vss out drv4 sky130_fd_pr__nfet_g5v0d10v5_YSH3F7
Xsky130_fd_pr__nfet_g5v0d10v5_YSH3F7_1 drv4 drv4 vss vss drv4 drv4 out vss drv4 drv4
+ vss drv4 out vss drv4 out vss out drv4 vss out drv4 sky130_fd_pr__nfet_g5v0d10v5_YSH3F7
Xsky130_fd_pr__nfet_g5v0d10v5_QCNVDG_0 vss crosscon vss crosscon drv4 drv4 vss drv4
+ crosscon crosscon crosscon vss sky130_fd_pr__nfet_g5v0d10v5_QCNVDG
Xsky130_fd_pr__pfet_g5v0d10v5_WECJAU_0 drv2 vdd_hi vdd_hi crosscon crosscon drv2 drv2
+ vdd_hi drv2 vdd_hi sky130_fd_pr__pfet_g5v0d10v5_WECJAU
Xsky130_fd_pr__pfet_g5v0d10v5_54K6JW_0 vdd_hi out out vdd_hi drv4 out drv4 vdd_hi
+ out vdd_hi drv4 drv4 drv4 vdd_hi drv4 out drv4 vdd_hi out drv4 vdd_hi out vdd_hi
+ drv4 drv4 drv4 vdd_hi drv4 drv4 out drv4 vdd_hi drv4 drv4 out vdd_hi out drv4 drv4
+ vdd_hi vdd_hi drv4 drv4 sky130_fd_pr__pfet_g5v0d10v5_54K6JW
Xsky130_fd_pr__pfet_g5v0d10v5_54K6JW_1 vdd_hi out out vdd_hi drv4 out drv4 vdd_hi
+ out vdd_hi drv4 drv4 drv4 vdd_hi drv4 out drv4 vdd_hi out drv4 vdd_hi out vdd_hi
+ drv4 drv4 drv4 vdd_hi drv4 drv4 out drv4 vdd_hi drv4 drv4 out vdd_hi out drv4 drv4
+ vdd_hi vdd_hi drv4 drv4 sky130_fd_pr__pfet_g5v0d10v5_54K6JW
Xsky130_fd_pr__pfet_g5v0d10v5_HKUKAU_0 in vdd_hi vdd_hi in drv1 drv1 sky130_fd_pr__pfet_g5v0d10v5_HKUKAU
Xsky130_fd_pr__pfet_g5v0d10v5_3QQKN5_1 vdd_hi vdd_hi drv2 vdd_hi drv1 drv1 sky130_fd_pr__pfet_g5v0d10v5_3QQKN5
.ends

.subckt sky130_fd_pr__nfet_01v8_U85QGS a_62_n200# a_n368_222# a_n224_n200# a_n320_n200#
+ a_398_222# a_n32_n200# a_n508_n200# a_302_n288# a_14_222# a_n464_n288# a_446_n200#
+ a_206_222# a_158_n200# a_110_n288# a_n272_n288# a_254_n200# a_n610_n374# a_n176_222#
+ a_350_n200# a_n416_n200# a_n128_n200# a_n80_n288#
X0 a_n128_n200# a_n176_222# a_n224_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1 a_n416_n200# a_n464_n288# a_n508_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2 a_n320_n200# a_n368_222# a_n416_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3 a_n32_n200# a_n80_n288# a_n128_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.32 pd=2.32 as=0.33 ps=2.33 w=2 l=0.15
X4 a_350_n200# a_302_n288# a_254_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5 a_254_n200# a_206_222# a_158_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6 a_158_n200# a_110_n288# a_62_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7 a_n224_n200# a_n272_n288# a_n320_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X8 a_446_n200# a_398_222# a_350_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X9 a_62_n200# a_14_222# a_n32_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.32 ps=2.32 w=2 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_B24TY6 a_n50_n298# a_50_n200# a_n108_n200# a_n266_n200#
+ w_n624_n496# a_n424_n200# a_108_n298# a_n208_n298# a_266_n298# a_208_n200# a_n366_n298#
+ a_366_n200#
X0 a_n108_n200# a_n208_n298# a_n266_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_208_n200# a_108_n298# a_50_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n266_n200# a_n366_n298# a_n424_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_366_n200# a_266_n298# a_208_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X4 a_50_n200# a_n50_n298# a_n108_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_ARHMTT a_n148_n1000# a_n386_n1000# a_566_n1000#
+ a_328_n1000# a_90_n1000# a_n758_n1222# a_n566_n1088# a_n328_n1088# a_n624_n1000#
+ a_n90_n1088# a_386_n1088# a_148_n1088#
X0 a_n148_n1000# a_n328_n1088# a_n386_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X1 a_90_n1000# a_n90_n1088# a_n148_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X2 a_566_n1000# a_386_n1088# a_328_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.9
X3 a_328_n1000# a_148_n1088# a_90_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X4 a_n386_n1000# a_n566_n1088# a_n624_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.9
.ends

.subckt audiodac_drv_ls in_p in_n out_p out_n vdd_hi vdd_lo VSUBS
XXM1 VSUBS in_p a_n3307_n18881# VSUBS in_p a_n3307_n18881# VSUBS in_p in_p in_p VSUBS
+ in_p a_n3307_n18881# in_p in_p VSUBS VSUBS in_p a_n3307_n18881# a_n3307_n18881#
+ VSUBS in_p sky130_fd_pr__nfet_01v8_U85QGS
XXM5 out_n vdd_hi out_p vdd_hi vdd_hi out_p out_n out_n out_n out_p out_n vdd_hi sky130_fd_pr__pfet_g5v0d10v5_B24TY6
XXM6 out_p vdd_hi out_n vdd_hi vdd_hi out_n out_p out_p out_p out_n out_p vdd_hi sky130_fd_pr__pfet_g5v0d10v5_B24TY6
Xsky130_fd_pr__nfet_05v0_nvt_ARHMTT_0 out_n a_n3307_n18881# a_n3307_n18881# out_n
+ a_n3307_n18881# VSUBS vdd_lo vdd_lo out_n vdd_lo vdd_lo vdd_lo sky130_fd_pr__nfet_05v0_nvt_ARHMTT
Xsky130_fd_pr__nfet_01v8_U85QGS_0 VSUBS in_n m1_n1994_n18882# VSUBS in_n m1_n1994_n18882#
+ VSUBS in_n in_n in_n VSUBS in_n m1_n1994_n18882# in_n in_n VSUBS VSUBS in_n m1_n1994_n18882#
+ m1_n1994_n18882# VSUBS in_n sky130_fd_pr__nfet_01v8_U85QGS
Xsky130_fd_pr__nfet_05v0_nvt_ARHMTT_1 m1_n1994_n18882# out_p out_p m1_n1994_n18882#
+ out_p VSUBS vdd_lo vdd_lo m1_n1994_n18882# vdd_lo vdd_lo vdd_lo sky130_fd_pr__nfet_05v0_nvt_ARHMTT
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VDASXE a_n1058_n5500# a_n1000_n5597# w_n1258_n5797#
+ a_1000_n5500#
X0 a_1000_n5500# a_n1000_n5597# a_n1058_n5500# w_n1258_n5797# sky130_fd_pr__pfet_g5v0d10v5 ad=15.95 pd=110.58 as=15.95 ps=110.58 w=55 l=10
.ends

.subckt sky130_iic_ip__audiodac_drv_lite in_p in_n out_p out_n in_hi vdd vss
Xaudiodac_drv_latch_0 audiodac_drv_latch_0/in_p audiodac_drv_latch_0/in_n vdd vss
+ audiodac_drv_latch
Xaudiodac_drv_lite_half_0 audiodac_drv_ls_0/out_n audiodac_drv_latch_0/in_n out_n
+ vdd vss audiodac_drv_lite_half
Xaudiodac_drv_lite_half_1 audiodac_drv_ls_0/out_p audiodac_drv_latch_0/in_p out_p
+ vdd vss audiodac_drv_lite_half
Xaudiodac_drv_ls_0 in_p in_n audiodac_drv_ls_0/out_p audiodac_drv_ls_0/out_n vdd in_hi
+ vss audiodac_drv_ls
Xsky130_fd_pr__pfet_g5v0d10v5_VDASXE_0 vdd vss vdd vdd sky130_fd_pr__pfet_g5v0d10v5_VDASXE
Xsky130_fd_pr__pfet_g5v0d10v5_VDASXE_1 vdd vss vdd vdd sky130_fd_pr__pfet_g5v0d10v5_VDASXE
.ends

.subckt comparator_bias VBN VSS VDD VBP ena3v3
X0 a_508213_646247# a_512471_646247# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X1 a_508213_647837# a_512471_648367# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X2 a_508215_648897# a_512471_648367# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X3 VSS VSS VBP VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X4 a_508215_648897# VDD VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X5 a_508213_647837# a_512471_647307# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X6 VSS VSS a_513709_648116# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X7 VDD VBP VBP VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X8 a_508213_646777# a_512471_646247# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X9 a_513709_648116# a_508213_646247# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X10 VBP VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X11 a_514109_648213# a_513709_648116# a_508213_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X12 a_513709_648116# a_508213_646247# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X13 a_514109_648213# a_513709_648116# a_508213_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X14 VSS VBN VBN VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X15 VDD a_508213_646247# a_513709_648116# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X16 VDD a_508213_646247# a_513709_648116# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X17 a_508213_646777# a_512471_647307# VDD sky130_fd_pr__res_high_po_1p41 l=19.29
X18 a_508213_646247# a_513709_648116# a_514109_648213# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X19 a_508213_646247# a_513709_648116# a_514109_648213# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X20 VBN ena3v3 a_514109_648213# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X21 a_513709_648116# VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X22 VBN VBN a_508213_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_58RHGH a_n108_n50# a_50_n50# a_n50_n147# w_n308_n347#
X0 a_50_n50# a_n50_n147# a_n108_n50# w_n308_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_99SHXG a_n1345_n531# a_629_n531# a_n629_n557#
+ a_n2003_n531# a_687_n557# a_n1287_n557# a_n29_n531# a_1287_n531# a_1345_n557# a_n687_n531#
+ a_n1945_n557# a_29_n557# a_1945_n531# VSUBS
X0 a_629_n531# a_29_n557# a_n29_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X1 a_n29_n531# a_n629_n557# a_n687_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X2 a_n1345_n531# a_n1945_n557# a_n2003_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=3
X3 a_n687_n531# a_n1287_n557# a_n1345_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X4 a_1945_n531# a_1345_n557# a_1287_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=3
X5 a_1287_n531# a_687_n557# a_629_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HHDTQV a_1945_n464# a_1345_n561# a_n1345_n464#
+ w_n2039_n564# a_629_n464# a_n1945_n561# a_29_n561# a_n2003_n464# a_n29_n464# a_1287_n464#
+ a_n629_n561# a_687_n561# a_n1287_n561# a_n687_n464#
X0 a_1287_n464# a_687_n561# a_629_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X1 a_1945_n464# a_1345_n561# a_1287_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=3
X2 a_629_n464# a_29_n561# a_n29_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X3 a_n29_n464# a_n629_n561# a_n687_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X4 a_n1345_n464# a_n1945_n561# a_n2003_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=3
X5 a_n687_n464# a_n1287_n561# a_n1345_n464# w_n2039_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H9Q64V a_n945_n531# a_n487_n531# a_n1345_n557#
+ a_1345_n531# a_n29_n531# a_887_n531# a_n887_n557# a_429_n531# a_945_n557# a_n429_n557#
+ a_487_n557# a_29_n557# a_n1403_n531# VSUBS
X0 a_429_n531# a_29_n557# a_n29_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1 a_887_n531# a_487_n557# a_429_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_n487_n531# a_n887_n557# a_n945_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X3 a_n29_n531# a_n429_n557# a_n487_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 a_1345_n531# a_945_n557# a_887_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X5 a_n945_n531# a_n1345_n557# a_n1403_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_SK4LJA a_n800_n561# a_800_n464# w_n894_n564#
+ a_n858_n464#
X0 a_800_n464# a_n800_n561# a_n858_n464# w_n894_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VKQJ4Z a_n1403_n464# a_945_n561# a_n429_n561#
+ a_487_n561# a_n945_n464# a_29_n561# a_n487_n464# a_1345_n464# a_n29_n464# a_887_n464#
+ a_429_n464# a_n1345_n561# w_n1439_n564# a_n887_n561#
X0 a_1345_n464# a_945_n561# a_887_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1 a_n945_n464# a_n1345_n561# a_n1403_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X2 a_429_n464# a_29_n561# a_n29_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X3 a_887_n464# a_487_n561# a_429_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 a_n487_n464# a_n887_n561# a_n945_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X5 a_n29_n464# a_n429_n561# a_n487_n464# w_n1439_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CNFY23 a_800_n531# a_n800_n557# a_n858_n531#
+ VSUBS
X0 a_800_n531# a_n800_n557# a_n858_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FXMKC5 a_n437_n531# a_n29_n531# a_379_n531# a_n379_n557#
+ a_29_n557# VSUBS
X0 a_379_n531# a_29_n557# a_n29_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1.75
X1 a_n29_n531# a_n379_n557# a_n437_n531# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1.75
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_H998DU a_129_n964# a_29_n1061# w_n223_n1064#
+ a_n129_n1061# a_n29_n964# a_n187_n964#
X0 a_n29_n964# a_n129_n1061# a_n187_n964# w_n223_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X1 a_129_n964# a_29_n1061# a_n29_n964# w_n223_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt comparator_core_cload VOUT DVDD VBN VSS VDD VINM VINP VBP CLOAD ena3v3
Xsky130_fd_pr__pfet_g5v0d10v5_58RHGH_0 VDD voutanalog ena3v3 VDD sky130_fd_pr__pfet_g5v0d10v5_58RHGH
Xsky130_fd_pr__nfet_g5v0d10v5_99SHXG_0 m3_516006_639184# VSS a_512694_640217# VSS
+ a_512694_640217# a_512694_640217# m3_516006_639184# m3_516006_639184# a_512694_640217#
+ VSS a_512694_640217# a_512694_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_99SHXG
Xsky130_fd_pr__pfet_g5v0d10v5_HHDTQV_0 VDD a_512178_641405# voutanalog VDD VDD a_512178_641405#
+ a_512178_641405# VDD voutanalog voutanalog a_512178_641405# a_512178_641405# a_512178_641405#
+ VDD sky130_fd_pr__pfet_g5v0d10v5_HHDTQV
Xsky130_fd_pr__nfet_g5v0d10v5_H9Q64V_0 voutanalog VSS a_512178_643337# VSS voutanalog
+ voutanalog a_512178_643337# VSS a_512178_643337# a_512178_643337# a_512178_643337#
+ a_512178_643337# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_H9Q64V
Xsky130_fd_pr__pfet_g5v0d10v5_SK4LJA_0 VBN a_508972_643337# VDD a_509888_643337# sky130_fd_pr__pfet_g5v0d10v5_SK4LJA
Xsky130_fd_pr__pfet_g5v0d10v5_SK4LJA_1 VBN a_509888_643337# VDD a_508972_643337# sky130_fd_pr__pfet_g5v0d10v5_SK4LJA
Xsky130_fd_pr__pfet_g5v0d10v5_VKQJ4Z_0 VDD a_509430_640243# a_509430_640243# a_509430_640243#
+ voutanalog a_509430_640243# VDD VDD voutanalog voutanalog VDD a_509430_640243# VDD
+ a_509430_640243# sky130_fd_pr__pfet_g5v0d10v5_VKQJ4Z
Xsky130_fd_pr__nfet_g5v0d10v5_CNFY23_0 a_508972_641405# VBP a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5_CNFY23
Xsky130_fd_pr__nfet_g5v0d10v5_FXMKC5_0 voutanalog m3_516006_639184# voutanalog VBP
+ VBP VSS sky130_fd_pr__nfet_g5v0d10v5_FXMKC5
Xsky130_fd_pr__pfet_g5v0d10v5_H998DU_0 VDD voutanalog VDD voutanalog a_515760_641405#
+ VDD sky130_fd_pr__pfet_g5v0d10v5_H998DU
Xsky130_fd_pr__nfet_g5v0d10v5_CNFY23_1 a_509888_641405# VBP a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5_CNFY23
X0 VSS CLOAD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X2 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X3 VOUT a_515760_641405# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X4 a_508572_644406# a_508572_644406# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X5 VOUT a_515760_641405# DVDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=3.1 ps=20.62 w=10 l=2
X6 a_508572_644406# VINM a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X7 VSS a_509030_640217# a_509430_640243# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X8 VSS a_512694_640217# a_512694_640217# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=5.58 w=5 l=3
X9 a_509030_640217# VINM a_509888_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X10 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X11 a_512694_640217# a_512694_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=5.58 as=0.725 ps=5.29 w=5 l=3
X12 VDD CLOAD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X13 VDD CLOAD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X14 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X15 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X16 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X17 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X18 VDD VDD a_509888_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X19 VSS VSS a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X20 VDD a_508572_644406# a_512694_640217# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=5.58 w=5 l=3
X21 a_512178_641405# a_512178_641405# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X22 a_509888_641405# VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X23 a_509888_643337# VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X24 a_512178_641405# VINP a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X25 a_512178_643337# VINP a_509888_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X26 a_512178_641405# VINP a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X27 a_512178_643337# VINP a_509888_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X28 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X29 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X30 a_512178_643337# a_512178_643337# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X31 VDD a_512178_641405# a_512178_641405# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X32 a_509888_643337# VINP a_512178_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X33 a_509888_641405# VINP a_512178_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X34 a_509888_641405# VINP a_512178_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X35 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=2
X36 VSS CLOAD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X37 a_509888_643337# VINP a_512178_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X38 a_509430_640243# a_509030_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X39 VSS a_509030_640217# a_509030_640217# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X40 a_512694_640217# a_508572_644406# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=5.58 as=0.725 ps=5.29 w=5 l=3
X41 VSS a_512178_643337# a_512178_643337# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X42 a_509430_640243# a_509430_640243# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X43 a_508972_641405# VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X44 a_508972_643337# VBP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X45 a_509030_640217# VINM a_509888_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X46 a_508572_644406# VINM a_509888_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X47 VSS CLOAD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X48 VSS voutanalog a_515760_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X49 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=2
X50 VDD CLOAD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X51 VDD a_508572_644406# a_508572_644406# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X52 VDD a_509430_640243# a_509430_640243# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X53 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=2
X54 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X55 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=2
X56 VSS VBN a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X57 a_509888_641405# VINM a_508572_644406# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X58 VSS CLOAD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X59 a_509030_640217# a_509030_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X60 VDD VBP a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X61 a_509888_643337# VINM a_509030_640217# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X62 a_509888_641405# VINM a_508572_644406# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X63 VDD CLOAD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X64 a_509888_643337# VINM a_509030_640217# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_ef_ip__ccomp3v_cl VINM VINP VDD VSS DVDD VOUT CLOAD ENA DVSS
Xcomparator_bias_0 comparator_bias_0/VBN VSS VDD comparator_bias_0/VBP comparator_bias_0/ena3v3
+ comparator_bias
Xcomparator_core_cload_0 VOUT DVDD comparator_bias_0/VBN VSS VDD VINM VINP comparator_bias_0/VBP
+ CLOAD comparator_bias_0/ena3v3 comparator_core_cload
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 ENA DVDD DVSS VDD VDD comparator_bias_0/ena3v3 VDD
+ DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 ENA DVSS DVSS VDD VDD sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_0 DVSS DVSS VDD VDD sky130_fd_sc_hvl__decap_4
.ends

* Black-box entry subcircuit for sky130_aa_ip__programmable_pll abstract view
.subckt sky130_aa_ip__programmable_pll S6 UP_INPUT DN_INPUT S2 S3 UP_OUT DN_OUT ITAIL
+ S4 VCTRL_IN LF_OFFCHIP S5 OUT_CORE OUT_USB D12 D13 D14 D15 F_IN D0 D1 D2 D3 D4 D5
+ D6 D7 D8 D9 D10 D16 D17 D18 D19 OUTB OUT PRE_SCALAR S1 S7 DIV_OUT VDD VSS
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0 a_n252_n322# a_50_n100# a_n108_n100#
+ a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VHBZVD a_n400_n197# a_400_n100# w_n658_n397#
+ a_n458_n100#
X0 a_400_n100# a_n400_n197# a_n458_n100# w_n658_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLNSY6 a_n29_n100# w_n387_n397# a_n187_n100#
+ a_29_n197# a_n129_n197# a_129_n100#
X0 a_129_n100# a_29_n197# a_n29_n100# w_n387_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n197# a_n187_n100# w_n387_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0 a_50_n400# a_n247_n622# a_n108_n400#
+ a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n247_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6 a_n50_n297# a_50_n200# w_n308_n497# a_n108_n200#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n308_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt mux2to1 A1 A0 Z VCC S VSS
XXM12 VSS m2_844_n775# VSS S sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM13 S m2_844_n775# VCC VCC sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6
XXM1 S Z VCC A0 sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6
XXM2 VSS Z A0 m2_844_n775# sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM3 m2_844_n775# Z VCC A1 sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6
XXM4 VSS Z A1 S sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YYAQG7 a_100_n200# a_n292_n422# a_n158_n200#
+ a_n100_n288#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n292_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0 a_n50_n197# a_50_n100# w_n308_n397#
+ a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T4TNG7 a_n100_n597# a_n100_21# a_100_109# a_100_n509#
+ a_n158_n509# a_n158_109# a_n297_n731#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n297_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n297_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_SALWK2 a_n88_n400# a_n33_n488# a_n190_n574# a_30_n400#
X0 a_30_n400# a_n33_n488# a_n88_n400# a_n190_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_FVGVKR a_n284_684# a_214_n1116# a_n118_684#
+ a_48_n1116# a_n284_n1116# a_n414_n1246# a_n118_n1116# a_48_684# a_214_684#
X0 a_214_684# a_214_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X1 a_n284_684# a_n284_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X2 a_48_684# a_48_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X3 a_n118_684# a_n118_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KL3SY6 a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_KB5CJD m3_n1186_n1040# c1_n1146_n1000#
X0 c1_n1146_n1000# m3_n1186_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__nfet_01v8_B8TQK3 a_n100_n597# a_n100_21# a_n260_n683# a_100_109#
+ a_100_n509# a_n158_n509# a_n158_109#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n260_n683# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n260_n683# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt comparator_final Vinn Vinp RST AVDD DVDD VSS
XXM12 VSS m2_9611_n3541# VSS vo1 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM23 m2_26_n3922# m2_26_n3922# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM13 m2_9611_n3541# AVDD AVDD vo1 vo1 AVDD sky130_fd_pr__pfet_g5v0d10v5_KLNSY6
XXM14 vo1 VSS VSS vo sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0
Xx1 VD VS VY AVDD vo1 VSS mux2to1
XXM25 VSS VSS vbn vbn sky130_fd_pr__nfet_g5v0d10v5_YYAQG7
XXM24 m2_26_n3922# vbn AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM15 vo vo1 li_9669_n4446# li_9669_n4446# sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM26 vbn vbn m2_1724_n5235# m2_1724_n5235# m2_26_n3922# m2_26_n3922# VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM16 VSS RST VSS m2_9611_n3541# sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM27 m2_26_n3922# VSS vbn m2_n888_n4722# sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0
XXM17 RST DVDD DVDD m2_9611_n3541# m2_9611_n3541# DVDD sky130_fd_pr__pfet_g5v0d10v5_KLNSY6
XXM28 VSS vbn VSS m2_n888_n4722# sky130_fd_pr__nfet_01v8_SALWK2
XXM19 li_9669_n4446# li_9669_n4446# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXR12 m1_2193_n3581# VSS m1_2193_n3581# m1_2360_n5380# m2_1724_n5235# VSS m1_2360_n5380#
+ m1_2525_n3581# m1_2525_n3581# sky130_fd_pr__res_xhigh_po_0p35_FVGVKR
XXM1 vbn vbn VS VS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM2 m1_7183_n5366# vt AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_1 vt vo sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM3 m1_7183_n5366# m1_7183_n5366# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
XXM4 m1_7183_n5366# VSS m2_6521_n3805# AVDD sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0
XXM5 m1_n1718_n3574# m1_n1718_n3574# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM6 vbn vbn VSS VSS vo vo VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM7 vt AVDD AVDD vo sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
XXM8 vt VSS VD AVDD sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0
Xsky130_fd_pr__nfet_01v8_B8TQK3_0 Vinn Vinn VSS VY VY VD VD sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_01v8_B8TQK3_1 Vinn Vinn VSS VS VS VD VD sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_01v8_B8TQK3_2 Vinn Vinn VSS VS VY VD VD sky130_fd_pr__nfet_01v8_B8TQK3
XXM20 m2_n888_n4722# m2_n888_n4722# AVDD m1_n1844_n4683# sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM10 Vinp Vinp VSS m2_6521_n3805# m2_6521_n3805# VS VS sky130_fd_pr__nfet_01v8_B8TQK3
XXM11 m1_n1844_n4683# m1_n1718_n3574# AVDD m1_n1844_n4683# sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n224# a_n73_n50# a_n33_n154# a_15_n50#
X0 a_15_n50# a_n33_n154# a_n73_n50# a_n175_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XPC8Y6 a_n29_n100# a_n187_n100# a_29_n197# a_n129_n197#
+ a_129_n100# w_n325_n319#
X0 a_129_n100# a_29_n197# a_n29_n100# w_n325_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n197# a_n187_n100# w_n325_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_GHZ9W9 a_n29_n100# a_89_n100# a_26_n197# w_n285_n319#
+ a_n92_n197# a_n147_n100#
X0 a_n29_n100# a_n92_n197# a_n147_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1 a_89_n100# a_26_n197# a_n29_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_2V27AY m4_200_n17880# c2_280_n17800# c2_n4018_n17800#
+ m4_n4098_n17880#
X0 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X1 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X2 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X3 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X4 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X5 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X6 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X7 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X8 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X9 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X10 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X11 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X12 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X13 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X14 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X15 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X16 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X17 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X18 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X19 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
.ends

.subckt sky130_fd_pr__nfet_01v8_PR763Z a_591_n50# a_1071_n50# a_207_n50# a_n465_n50#
+ a_n207_n76# a_n945_n50# a_783_n50# a_1263_n50# a_n177_n50# a_n1299_72# a_n1427_n224#
+ a_n657_n50# a_n1137_n50# a_n1325_n50# a_495_n50# a_111_n50# a_975_n50# a_n369_n50#
+ a_n975_n76# a_n849_n50# a_1167_n50# a_687_n50# a_303_n50# a_n561_n50# a_n1041_n50#
+ a_n1167_n76# a_n81_n50# a_399_n50# a_879_n50# a_n273_n50# a_15_n50# a_n753_n50#
+ a_n1233_n50#
X0 a_15_n50# a_n207_n76# a_n81_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X1 a_111_n50# a_n207_n76# a_15_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X2 a_n273_n50# a_n975_n76# a_n369_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X3 a_n81_n50# a_n207_n76# a_n177_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X4 a_n177_n50# a_n207_n76# a_n273_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X5 a_303_n50# a_n207_n76# a_207_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X6 a_591_n50# a_n207_n76# a_495_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X7 a_207_n50# a_n207_n76# a_111_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X8 a_399_n50# a_n207_n76# a_303_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X9 a_495_n50# a_n207_n76# a_399_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X10 a_687_n50# a_n207_n76# a_591_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X11 a_783_n50# a_n207_n76# a_687_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X12 a_975_n50# a_n207_n76# a_879_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X13 a_n1041_n50# a_n1167_n76# a_n1137_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X14 a_879_n50# a_n207_n76# a_783_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X15 a_n1233_n50# a_n1299_72# a_n1325_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X16 a_n1137_n50# a_n1167_n76# a_n1233_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X17 a_n561_n50# a_n975_n76# a_n657_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X18 a_1071_n50# a_n207_n76# a_975_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X19 a_1167_n50# a_n207_n76# a_1071_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X20 a_1263_n50# a_n207_n76# a_1167_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X21 a_n945_n50# a_n975_n76# a_n1041_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X22 a_n849_n50# a_n975_n76# a_n945_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X23 a_n753_n50# a_n975_n76# a_n849_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X24 a_n657_n50# a_n975_n76# a_n753_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X25 a_n465_n50# a_n975_n76# a_n561_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X26 a_n369_n50# a_n975_n76# a_n465_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_DD63S8 a_n465_n202# a_n945_18# a_1167_n202# a_n81_18#
+ a_n273_18# a_15_n202# a_n561_n202# a_975_18# a_n177_n202# a_303_18# a_1263_n202#
+ a_879_n202# a_111_n202# a_n1041_18# a_n975_n299# a_n273_n202# a_n1137_n202# a_n849_18#
+ a_975_n202# a_n561_18# a_1071_18# a_879_18# a_n177_18# a_n1233_n202# a_207_18# a_591_18#
+ a_1071_n202# a_687_n202# a_15_18# a_n465_18# a_783_n202# a_399_n202# a_n81_n202#
+ a_n849_n202# w_n1463_n397# a_495_18# a_n1233_18# a_n1041_n202# a_n1299_n299# a_495_n202#
+ a_n945_n202# a_n753_18# a_1263_18# a_n369_18# a_783_18# a_n1137_18# a_n207_n299#
+ a_591_n202# a_n657_n202# a_399_18# a_111_18# a_207_n202# a_n1167_n299# a_n753_n202#
+ a_n1325_n202# a_1167_18# a_n657_18# a_n369_n202# a_n1325_18# a_303_n202# a_687_18#
X0 a_n1233_n202# a_n1299_n299# a_n1325_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_591_n202# a_n207_n299# a_495_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X2 a_n657_18# a_n975_n299# a_n753_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X3 a_975_18# a_n207_n299# a_879_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X4 a_1263_18# a_n207_n299# a_1167_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X5 a_n849_n202# a_n975_n299# a_n945_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X6 a_n945_18# a_n975_n299# a_n1041_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X7 a_879_18# a_n207_n299# a_783_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X8 a_n177_n202# a_n207_n299# a_n273_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X9 a_207_n202# a_n207_n299# a_111_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X10 a_1167_18# a_n207_n299# a_1071_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X11 a_n1137_n202# a_n1167_n299# a_n1233_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X12 a_495_n202# a_n207_n299# a_399_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X13 a_n849_18# a_n975_n299# a_n945_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X14 a_n81_18# a_n207_n299# a_n177_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X15 a_n561_n202# a_n975_n299# a_n657_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X16 a_111_n202# a_n207_n299# a_15_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X17 a_783_n202# a_n207_n299# a_687_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X18 a_1071_n202# a_n207_n299# a_975_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X19 a_303_18# a_n207_n299# a_207_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X20 a_399_n202# a_n207_n299# a_303_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X21 a_n1041_18# a_n1167_n299# a_n1137_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X22 a_n273_18# a_n975_n299# a_n369_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X23 a_111_18# a_n207_n299# a_15_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X24 a_n465_n202# a_n975_n299# a_n561_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X25 a_687_n202# a_n207_n299# a_591_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X26 a_207_18# a_n207_n299# a_111_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X27 a_591_18# a_n207_n299# a_495_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X28 a_n753_n202# a_n975_n299# a_n849_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X29 a_975_n202# a_n207_n299# a_879_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X30 a_n177_18# a_n207_n299# a_n273_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X31 a_15_18# a_n207_n299# a_n81_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X32 a_n81_n202# a_n207_n299# a_n177_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X33 a_1263_n202# a_n207_n299# a_1167_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X34 a_n561_18# a_n975_n299# a_n657_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X35 a_495_18# a_n207_n299# a_399_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X36 a_15_n202# a_n207_n299# a_n81_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X37 a_n1233_18# a_n1299_n299# a_n1325_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X38 a_n1041_n202# a_n1167_n299# a_n1137_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X39 a_n369_n202# a_n975_n299# a_n465_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X40 a_n465_18# a_n975_n299# a_n561_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X41 a_399_18# a_n207_n299# a_303_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X42 a_n657_n202# a_n975_n299# a_n753_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X43 a_n1137_18# a_n1167_n299# a_n1233_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X44 a_783_18# a_n207_n299# a_687_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X45 a_879_n202# a_n207_n299# a_783_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X46 a_1071_18# a_n207_n299# a_975_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X47 a_n945_n202# a_n975_n299# a_n1041_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X48 a_1167_n202# a_n207_n299# a_1071_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X49 a_n753_18# a_n975_n299# a_n849_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X50 a_n369_18# a_n975_n299# a_n465_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X51 a_303_n202# a_n207_n299# a_207_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X52 a_687_18# a_n207_n299# a_591_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X53 a_n273_n202# a_n975_n299# a_n369_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt por_output_buffer w_33421_n285686# m2_34641_n286220# VSUBS m1_33354_n286009#
XXM53 m2_34641_n286220# VSUBS m2_34641_n286220# VSUBS m2_33873_n286220# m2_33873_n286220#
+ m2_34641_n286220# VSUBS m2_34641_n286220# m1_33354_n286009# VSUBS VSUBS m2_33681_n286220#
+ m2_33489_n286220# VSUBS VSUBS m2_34641_n286220# m2_33873_n286220# m2_33681_n286220#
+ VSUBS m2_34641_n286220# VSUBS VSUBS m2_33873_n286220# VSUBS m2_33489_n286220# VSUBS
+ m2_34641_n286220# VSUBS VSUBS m2_34641_n286220# m2_33873_n286220# VSUBS sky130_fd_pr__nfet_01v8_PR763Z
XXM54 w_33421_n285686# m2_33873_n286220# m2_34641_n286220# w_33421_n285686# w_33421_n285686#
+ m2_34641_n286220# m2_33873_n286220# m2_34641_n286220# m2_34641_n286220# w_33421_n285686#
+ w_33421_n285686# w_33421_n285686# w_33421_n285686# w_33421_n285686# m2_33681_n286220#
+ w_33421_n285686# m2_33681_n286220# w_33421_n285686# m2_34641_n286220# m2_33873_n286220#
+ w_33421_n285686# w_33421_n285686# m2_34641_n286220# w_33421_n285686# m2_34641_n286220#
+ m2_34641_n286220# w_33421_n285686# w_33421_n285686# m2_34641_n286220# w_33421_n285686#
+ m2_34641_n286220# m2_34641_n286220# w_33421_n285686# w_33421_n285686# w_33421_n285686#
+ w_33421_n285686# w_33421_n285686# w_33421_n285686# m1_33354_n286009# w_33421_n285686#
+ m2_33873_n286220# m2_33873_n286220# w_33421_n285686# m2_33873_n286220# m2_34641_n286220#
+ m2_33681_n286220# m2_33873_n286220# m2_34641_n286220# w_33421_n285686# m2_34641_n286220#
+ w_33421_n285686# m2_34641_n286220# m2_33489_n286220# m2_33873_n286220# m2_33489_n286220#
+ m2_34641_n286220# w_33421_n285686# m2_33873_n286220# m2_33489_n286220# w_33421_n285686#
+ w_33421_n285686# sky130_fd_pr__pfet_01v8_DD63S8
.ends

.subckt sky130_fd_pr__pfet_01v8_U6B66J a_n73_118# a_n33_21# w_n211_n477# a_n73_n258#
+ a_15_118# a_n33_n355# a_15_n258#
X0 a_15_118# a_n33_21# a_n73_118# w_n211_n477# sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X1 a_15_n258# a_n33_n355# a_n73_n258# w_n211_n477# sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PQJ659 a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_01v8_G7LLWL a_n29_n50# a_26_n154# a_n249_n224# a_n147_n50#
+ a_89_n50# a_n92_n154#
X0 a_89_n50# a_26_n154# a_n29_n50# a_n249_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X1 a_n29_n50# a_n92_n154# a_n147_n50# a_n249_n224# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_5QNSAB a_n33_n50# a_n227_n224# a_63_n50# a_n125_n50#
+ a_n81_n154#
X0 a_n33_n50# a_n81_n154# a_n125_n50# a_n227_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X1 a_63_n50# a_n81_n154# a_n33_n50# a_n227_n224# sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLZS5A a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_01v8_SKYQWJ a_n88_n318# a_30_118# a_n33_n415# a_n33_21#
+ a_n88_118# a_30_n318# w_n226_n537#
X0 a_30_n318# a_n33_n415# a_n88_n318# w_n226_n537# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_30_118# a_n33_21# a_n88_118# w_n226_n537# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69TNYL a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSE8X6 a_n331_n402# a_29_n268# a_n29_n180# a_n129_n268#
+ a_n187_n180# a_129_n180#
X0 a_129_n180# a_29_n268# a_n29_n180# a_n331_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.5
X1 a_n29_n180# a_n129_n268# a_n187_n180# a_n331_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6 a_129_n290# a_29_n387# a_n129_n387# a_n29_n290#
+ a_n187_n290# w_n387_n587#
X0 a_129_n290# a_29_n387# a_n29_n290# w_n387_n587# sky130_fd_pr__pfet_g5v0d10v5 ad=0.841 pd=6.38 as=0.4205 ps=3.19 w=2.9 l=0.5
X1 a_n29_n290# a_n129_n387# a_n187_n290# w_n387_n587# sky130_fd_pr__pfet_g5v0d10v5 ad=0.4205 pd=3.19 as=0.841 ps=6.38 w=2.9 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_X6X8XQ a_n81_n167# a_n33_n70# a_63_n70# a_n125_n70#
+ w_n263_n289#
X0 a_n33_n70# a_n81_n167# a_n125_n70# w_n263_n289# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_63_n70# a_n81_n167# a_n33_n70# w_n263_n289# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N5F8XL a_n108_n180# a_n242_n402# a_n50_n268#
+ a_50_n180#
X0 a_50_n180# a_n50_n268# a_n108_n180# a_n242_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_FJFAMD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt levelShifter ain aout VCCL VCCH VSS
Xsky130_fd_pr__nfet_g5v0d10v5_WSE8X6_0 VSS S1B VSS S1B m2_2125_n529# m2_2125_n529#
+ sky130_fd_pr__nfet_g5v0d10v5_WSE8X6
XXM12 VSS S1 VSS S1 m1_2633_n381# m1_2633_n381# sky130_fd_pr__nfet_g5v0d10v5_WSE8X6
XXM13 m2_2125_n529# m1_2633_n381# m1_2633_n381# VCCH m2_2125_n529# VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
XXM1 ain VCCL S1 S1 VCCL sky130_fd_pr__pfet_01v8_X6X8XQ
XXM2 m1_2633_n381# m2_2125_n529# m2_2125_n529# VCCH m1_2633_n381# VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
XXM4 VSS VSS S1 S1B sky130_fd_pr__nfet_01v8_L9ESAD
XXM5 S1 VCCL S1B S1B VCCL sky130_fd_pr__pfet_01v8_X6X8XQ
XXM6 VSS VSS ain S1 sky130_fd_pr__nfet_01v8_L9ESAD
XXM7 aout VSS m2_2125_n529# VSS sky130_fd_pr__nfet_g5v0d10v5_N5F8XL
XXM8 aout m2_2125_n529# m2_2125_n529# VCCH aout VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
Xsky130_fd_pr__cap_mim_m3_1_FJFAMD_0 m2_2125_n529# VCCH sky130_fd_pr__cap_mim_m3_1_FJFAMD
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ESEQJ8 a_n282_n422# a_80_n200# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n282_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TBT74C c1_n1746_n1600# m3_n1786_n1640#
X0 c1_n1746_n1600# m3_n1786_n1640# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SYBQJL a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CAF9E7 a_29_n347# a_n129_n347# a_n29_n250# a_n187_n250#
+ w_n387_n547# a_129_n250#
X0 a_129_n250# a_29_n347# a_n29_n250# w_n387_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X1 a_n29_n250# a_n129_n347# a_n187_n250# w_n387_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_X6E435 a_n29_n100# a_n187_n100# a_129_n100# a_n331_n322#
+ a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n331_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n331_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X11 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X16 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X18 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X19 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X22 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X23 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X24 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X25 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X26 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X27 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X28 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X29 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X30 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X31 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt por_output_driver_h sky130_fd_sc_hvl__inv_16_0/VPWR sky130_fd_sc_hvl__inv_16_0/Y
+ sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_0/VGND sky130_fd_sc_hvl__inv_16_1/VPWR
+ m2_26866_n292108# m2_26862_n291518# sky130_fd_sc_hvl__inv_16_1/VGND sky130_fd_sc_hvl__inv_16_1/Y
+ VSUBS
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_0 m2_26960_n292468# m2_26960_n292468# m2_27646_n292468#
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_2 m2_27646_n292468# m2_27646_n292468# sky130_fd_sc_hvl__inv_16_1/A
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_1 m2_26866_n292108# m2_26866_n292108# m2_26960_n292468#
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_0 VSUBS m2_26960_n292468# m2_26960_n292468# VSUBS
+ m2_26866_n292108# m2_26866_n292108# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_2 VSUBS sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_1/A
+ VSUBS m2_27646_n292468# m2_27646_n292468# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_1 VSUBS m2_27646_n292468# m2_27646_n292468# VSUBS
+ m2_26960_n292468# m2_26960_n292468# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_sc_hvl__inv_16_0 sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_0/VGND
+ VSUBS sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_0/VPWR sky130_fd_sc_hvl__inv_16_0/Y
+ sky130_fd_sc_hvl__inv_16
Xsky130_fd_sc_hvl__inv_16_1 sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_1/VGND
+ VSUBS sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_1/VPWR sky130_fd_sc_hvl__inv_16_1/Y
+ sky130_fd_sc_hvl__inv_16
.ends

.subckt sky130_fd_pr__pfet_01v8_X6XW7S a_63_n258# a_n33_118# a_63_118# a_n125_118#
+ a_n33_n258# a_n81_21# w_n263_n477# a_n125_n258# a_n81_n355#
X0 a_n33_n258# a_n81_n355# a_n125_n258# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_n33_118# a_n81_21# a_n125_118# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X2 a_63_n258# a_n81_n355# a_n33_n258# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X3 a_63_118# a_n81_21# a_n33_118# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_RQPX7Z c2_n1869_n1600# m4_n1949_n1680#
X0 c2_n1869_n1600# m4_n1949_n1680# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_HYMU45 c2_n1069_n800# m4_n1149_n880#
X0 c2_n1069_n800# m4_n1149_n880# sky130_fd_pr__cap_mim_m3_2 l=8 w=8
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_4PHTN9 m4_n1349_n1080# c2_n1269_n1000#
X0 c2_n1269_n1000# m4_n1349_n1080# sky130_fd_pr__cap_mim_m3_2 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_EEU5EF m3_n4192_n17480# c1_n4152_n17440# c1_160_n17440#
+ m3_120_n17480#
X0 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X1 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X2 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X3 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X4 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X5 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X6 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X7 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X8 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X9 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X10 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X11 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X12 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X13 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X14 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X15 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X16 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X17 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X18 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X19 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_RRZ644 m3_n986_n840# c1_n946_n800#
X0 c1_n946_n800# m3_n986_n840# sky130_fd_pr__cap_mim_m3_1 l=8 w=8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_KA8C77 a_516_984# a_n2292_n1416# a_n1590_n1416#
+ a_2622_984# a_1218_n1416# a_n2760_n1416# a_282_n1416# a_n654_984# a_n888_984# a_48_n1416#
+ a_n420_984# a_n420_n1416# a_750_n1416# a_n2760_984# a_1686_984# a_1452_984# a_n2526_984#
+ a_1218_984# a_n2058_n1416# a_n1356_n1416# a_2388_n1416# a_1686_n1416# a_n1824_n1416#
+ a_n2526_n1416# a_n1590_984# a_n888_n1416# a_n2890_n1546# a_516_n1416# a_n1122_984#
+ a_n1356_984# a_282_984# a_2388_984# a_2154_984# a_1920_984# a_48_984# a_n1122_n1416#
+ a_2154_n1416# a_n186_n1416# a_n186_984# a_1452_n1416# a_2622_n1416# a_1920_n1416#
+ a_984_n1416# a_n654_n1416# a_n2292_984# a_984_984# a_n1824_984# a_750_984# a_n2058_984#
X0 a_n1590_984# a_n1590_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X1 a_282_984# a_282_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X2 a_1218_984# a_1218_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X3 a_2154_984# a_2154_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X4 a_n888_984# a_n888_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X5 a_1920_984# a_1920_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X6 a_750_984# a_750_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X7 a_2622_984# a_2622_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X8 a_n2760_984# a_n2760_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X9 a_516_984# a_516_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X10 a_n186_984# a_n186_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X11 a_n2292_984# a_n2292_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X12 a_n1356_984# a_n1356_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X13 a_n2058_984# a_n2058_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X14 a_1686_984# a_1686_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X15 a_n654_984# a_n654_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X16 a_n1824_984# a_n1824_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X17 a_2388_984# a_2388_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X18 a_n420_984# a_n420_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X19 a_n2526_984# a_n2526_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X20 a_984_984# a_984_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X21 a_n1122_984# a_n1122_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X22 a_48_984# a_48_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X23 a_1452_984# a_1452_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XSEQJ6 a_189_n200# a_407_n200# a_n599_n422# a_n189_n288#
+ a_29_n288# a_247_n288# a_n407_n288# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n288# a_n465_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X1 a_407_n200# a_247_n288# a_189_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_189_n200# a_29_n288# a_n29_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_n29_n200# a_n189_n288# a_n247_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_01v8_6QC8WZ a_n29_n100# a_89_n100# a_26_n197# w_n285_n319#
+ a_n92_n197# a_n147_n100#
X0 a_n29_n100# a_n92_n197# a_n147_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1 a_89_n100# a_26_n197# a_n29_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_sc_ls__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=1
.ends

.subckt sky130_fd_sc_ls__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 a_922_127# a_841_288# a_850_127# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_1598_93# a_1266_119# a_1736_119# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VGND a_1598_93# a_1550_119# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 a_33_74# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X4 a_1266_119# a_300_74# a_841_288# VNB sky130_fd_pr__nfet_01v8 ad=0.3067 pd=2.01 as=0.1073 ps=1.03 w=0.74 l=0.15
X5 a_1266_119# a_507_347# a_841_288# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22385 pd=1.7 as=0.39 ps=1.78 w=1 l=0.15
X6 a_714_127# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.07245 ps=0.765 w=0.42 l=0.15
X7 a_841_288# a_714_127# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.275 ps=2.55 w=1 l=0.15
X8 VPWR a_1266_119# a_1598_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0.063 ps=0.72 w=0.42 l=0.15
X9 a_714_127# a_507_347# a_33_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X10 a_507_347# a_300_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.40345 pd=2.86 as=0.295 ps=2.59 w=1 l=0.15
X11 VGND RESET_B a_120_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X12 VPWR a_1598_93# a_1547_508# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1550_119# a_507_347# a_1266_119# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.3067 ps=2.01 w=0.42 l=0.15
X14 a_1736_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X15 a_850_127# a_300_74# a_714_127# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X16 a_300_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2035 pd=2.03 as=0.1212 ps=1.1 w=0.74 l=0.15
X17 a_1547_508# a_300_74# a_1266_119# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.22385 ps=1.7 w=0.42 l=0.15
X18 a_1598_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_841_288# a_714_127# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1073 pd=1.03 as=0.240325 ps=1.715 w=0.74 l=0.15
X20 a_300_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.172775 ps=1.58 w=1 l=0.15
X21 VPWR a_841_288# a_817_463# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 a_120_74# D a_33_74# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X23 VPWR RESET_B a_33_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172775 pd=1.58 as=0.063 ps=0.72 w=0.42 l=0.15
X24 Q a_1934_94# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2146 pd=2.06 as=0.126075 ps=1.1 w=0.74 l=0.15
X25 a_817_463# a_507_347# a_714_127# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X26 VGND a_1266_119# a_1934_94# VNB sky130_fd_pr__nfet_01v8 ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X27 a_714_127# a_300_74# a_33_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X28 VGND RESET_B a_922_127# VNB sky130_fd_pr__nfet_01v8 ad=0.240325 pd=1.715 as=0.0441 ps=0.63 w=0.42 l=0.15
X29 a_507_347# a_300_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2479 pd=2.15 as=0.3299 ps=2.67 w=0.74 l=0.15
X30 VPWR a_1266_119# a_1934_94# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1862 pd=1.475 as=0.231 ps=2.23 w=0.84 l=0.15
X31 Q a_1934_94# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XJT6XQ a_n33_n50# a_63_n50# a_n125_n50# a_n81_n157#
+ w_n263_n269#
X0 a_n33_n50# a_n81_n157# a_n125_n50# w_n263_n269# sky130_fd_pr__pfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X1 a_63_n50# a_n81_n157# a_n33_n50# w_n263_n269# sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt TieH_1p8 TieH VSS VCC
XXM4 VSS m2_456_n646# m2_456_n646# VSS sky130_fd_pr__nfet_01v8_L9ESAD
XXM5 TieH VCC VCC m2_456_n646# VCC sky130_fd_pr__pfet_01v8_XJT6XQ
.ends

.subckt sky130_fd_sc_ls__buf_8 A VGND VNB VPB VPWR X
X0 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.2627 pd=2.19 as=0.10545 ps=1.025 w=0.74 l=0.15
X9 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X10 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X11 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X12 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1876 pd=1.455 as=0.168 ps=1.42 w=1.12 l=0.15
X15 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10545 pd=1.025 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X19 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
.ends

.subckt sky130_fd_sc_ls__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_30_78# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.05985 ps=0.705 w=0.42 l=0.15
X1 VGND RESET_B a_894_138# VNB sky130_fd_pr__nfet_01v8 ad=0.211225 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 a_894_138# a_830_359# a_816_138# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 VPWR a_1518_203# a_1468_493# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1864_409# a_1266_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5 a_830_359# a_695_457# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.24605 pd=1.405 as=0.211225 ps=1.45 w=0.74 l=0.15
X6 a_816_138# a_490_390# a_695_457# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X7 a_1476_81# a_306_96# a_1266_74# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X8 VGND a_1864_409# Q VNB sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_490_390# a_306_96# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.15 ps=1.3 w=1 l=0.15
X10 a_1468_493# a_490_390# a_1266_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X11 VPWR CLK a_306_96# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.31 ps=2.62 w=1 l=0.15
X12 a_1266_74# a_306_96# a_830_359# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23015 pd=1.73 as=0.190625 ps=1.505 w=1 l=0.15
X13 a_830_359# a_695_457# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.190625 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X14 VPWR a_1864_409# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X15 a_1656_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X16 VPWR a_1266_74# a_1518_203# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X17 a_1864_409# a_1266_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X18 VGND CLK a_306_96# VNB sky130_fd_pr__nfet_01v8 ad=0.162375 pd=1.255 as=0.2646 ps=2.4 w=0.74 l=0.15
X19 a_1518_203# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X20 a_695_457# a_306_96# a_30_78# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X21 a_1518_203# a_1266_74# a_1656_81# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_695_457# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1239 pd=1.43 as=0.137125 ps=1.155 w=0.42 l=0.15
X23 a_117_78# D a_30_78# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X24 VPWR a_830_359# a_785_457# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.137125 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X25 VGND a_1518_203# a_1476_81# VNB sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 VGND RESET_B a_117_78# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 a_785_457# a_306_96# a_695_457# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X28 a_695_457# a_490_390# a_30_78# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X29 a_30_78# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.1197 ps=1.41 w=0.42 l=0.15
X30 a_490_390# a_306_96# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2183 pd=2.07 as=0.162375 ps=1.255 w=0.74 l=0.15
X31 a_1266_74# a_490_390# a_830_359# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
.ends

.subckt sky130_fd_sc_ls__xor2_1 A B VGND VNB VPB VPWR X
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X4 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.177375 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.126075 ps=1.1 w=0.74 l=0.15
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8 ad=0.126075 pd=1.1 as=0.177375 ps=1.195 w=0.55 l=0.15
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8 ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
.ends

.subckt delayPulse_digital sky130_fd_sc_ls__dfrtp_1_0/RESET_B sky130_fd_sc_ls__dfrtp_1_0/CLK
+ sky130_fd_sc_ls__dfrtn_1_0/Q sky130_fd_sc_ls__dfrtp_1_0/Q sky130_fd_sc_ls__xor2_1_0/B
+ sky130_fd_sc_ls__xor2_1_0/A TieH_1p8_0/VCC VSUBS
Xsky130_fd_sc_ls__decap_4_0 VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__decap_4
Xsky130_fd_sc_ls__dfrtn_1_0 sky130_fd_sc_ls__buf_8_0/X TieH_1p8_0/TieH sky130_fd_sc_ls__dfrtp_1_0/CLK
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__dfrtn_1_0/Q sky130_fd_sc_ls__dfrtn_1
XTieH_1p8_0 TieH_1p8_0/TieH VSUBS TieH_1p8_0/VCC TieH_1p8
Xsky130_fd_sc_ls__buf_8_0 sky130_fd_sc_ls__buf_8_0/A VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC
+ sky130_fd_sc_ls__buf_8_0/X sky130_fd_sc_ls__buf_8
Xsky130_fd_sc_ls__dfrtp_1_0 sky130_fd_sc_ls__dfrtp_1_0/CLK TieH_1p8_0/TieH sky130_fd_sc_ls__dfrtp_1_0/RESET_B
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__dfrtp_1_0/Q sky130_fd_sc_ls__dfrtp_1
Xsky130_fd_sc_ls__xor2_1_0 sky130_fd_sc_ls__xor2_1_0/A sky130_fd_sc_ls__xor2_1_0/B
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__buf_8_0/A sky130_fd_sc_ls__xor2_1
.ends

.subckt delayPulse_final din por Vbg porb porb_h[0] porb_h[1] VCCH VCCL VSS
XXM34 VSS VSS m4_25183_n288425# m2_24504_n284758# sky130_fd_pr__nfet_01v8_L9ESAD
XXM23 m2_29747_n287456# m2_27024_n287466# vbp2 vbp2 m2_27024_n287466# VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM12 VT3 VCCL VT2 VCCL VT2 VCCL sky130_fd_pr__pfet_01v8_GHZ9W9
Xsky130_fd_pr__cap_mim_m3_2_2V27AY_0 VT3 VSS VSS VT3 sky130_fd_pr__cap_mim_m3_2_2V27AY
Xpor_output_buffer_1 VCCL por VSS porPre por_output_buffer
XXM35 VCCL m4_25183_n288425# VCCL VCCL m2_24504_n284758# m4_25183_n288425# m2_24504_n284758#
+ sky130_fd_pr__pfet_01v8_U6B66J
XXM24 m2_23680_n288167# m2_23680_n288167# VCCH m1_22999_n287228# sky130_fd_pr__pfet_g5v0d10v5_PQJ659
XXM13 m2_31224_n287586# VT3 VSS VSS VSS VT3 sky130_fd_pr__nfet_01v8_G7LLWL
Xsky130_fd_pr__cap_mim_m3_2_2V27AY_1 VT2 VSS VSS VT2 sky130_fd_pr__cap_mim_m3_2_2V27AY
XXM36 VSS VSS Td_Sd Td_Sd m2_24748_n284671# sky130_fd_pr__nfet_01v8_5QNSAB
XXM25 m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# VCCH
+ m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# VCCH m1_22999_n287228# m1_22999_n287228#
+ m1_22999_n287228# m1_22999_n287228# VCCH VCCH VCCH m1_22999_n287228# VCCH sky130_fd_pr__pfet_g5v0d10v5_KLZS5A
XXM14 m2_29747_n287456# m2_31224_n287586# VT3 VT3 m2_29747_n287456# m2_31224_n287586#
+ m2_29747_n287456# sky130_fd_pr__pfet_01v8_SKYQWJ
XXM26 m1_22125_n286949# VSS m2_23680_n288167# Vbg sky130_fd_pr__nfet_g5v0d10v5_69TNYL
Xx3 porbPre x3/aout VCCL VCCH VSS levelShifter
XXM38 VSS VSS m2_24504_n284758# m2_24748_n284671# sky130_fd_pr__nfet_01v8_L9ESAD
XXM27 VSS VSS m2_31224_n287586# m2_31884_n287663# sky130_fd_pr__nfet_01v8_L9ESAD
XXM16 m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM39 VCCL m2_24504_n284758# VCCL VCCL m2_24748_n284671# m2_24504_n284758# m2_24748_n284671#
+ sky130_fd_pr__pfet_01v8_U6B66J
XXM17 VSS vbp2 VSS vbn1 sky130_fd_pr__nfet_g5v0d10v5_ESEQJ8
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_0 vbp1 VCCL sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM29 VCCL m2_31224_n287586# VCCL VCCL m2_31884_n287663# m2_31224_n287586# m2_31884_n287663#
+ sky130_fd_pr__pfet_01v8_U6B66J
XXM18 m1_22999_n287228# VCCH VCCH m2_24152_n287606# sky130_fd_pr__pfet_g5v0d10v5_PQJ659
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_1 vbn1 VSS sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM19 vbn1 VSS vbn1 VSS VSS vbn1 vbn1 vbn1 vbn1 vbn1 vbn1 vbn1 VSS vbn1 VSS vbn1 sky130_fd_pr__nfet_g5v0d10v5_SYBQJL
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_2 m1_22999_n287228# VCCH sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM1 vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM2 VCCL m2_30306_n287752# din din VCCL m2_30306_n287752# VCCL sky130_fd_pr__pfet_01v8_SKYQWJ
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_0 VSS m4_25183_n288425# sky130_fd_pr__cap_mim_m3_1_KB5CJD
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_1 VSS m2_24748_n284671# sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM3 VCCL Td_S m2_30306_n287752# m2_30306_n287752# VCCL Td_S VCCL sky130_fd_pr__pfet_01v8_SKYQWJ
XXM4 Td_Lb VSS VSS VSS Td_L sky130_fd_pr__nfet_01v8_5QNSAB
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_2 VSS m2_24504_n284758# sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM5 VT2 m2_30306_n287752# VSS VSS VSS m2_30306_n287752# sky130_fd_pr__nfet_01v8_G7LLWL
XXM6 VT3 VT2 VSS m2_29342_n288187# m2_29342_n288187# VT2 sky130_fd_pr__nfet_01v8_G7LLWL
Xpor_output_driver_h_0 VCCH porb_h[0] VCCH VSS VCCH x3/aout VCCH VSS porb_h[1] VSS
+ por_output_driver_h
XXM7 VSS din VSS m2_30306_n287752# m2_30306_n287752# din sky130_fd_pr__nfet_01v8_G7LLWL
XXM8 VSS m2_30306_n287752# VSS Td_S Td_S m2_30306_n287752# sky130_fd_pr__nfet_01v8_G7LLWL
XXM9 VCCL Td_Lb VCCL VCCL Td_Lb Td_L VCCL VCCL Td_L sky130_fd_pr__pfet_01v8_X6XW7S
Xsky130_fd_pr__cap_mim_m3_2_RQPX7Z_0 VCCL vbp1 sky130_fd_pr__cap_mim_m3_2_RQPX7Z
XXC1 VSS vbn1 sky130_fd_pr__cap_mim_m3_2_RQPX7Z
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[0] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[1] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[2] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[3] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[4] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[5] VCCL m2_29064_n286804# vbp1 vbp1 m2_29064_n286804#
+ VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[6] m2_29759_n286901# m2_29064_n286804# vbp2 vbp2
+ m2_29064_n286804# VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXC3 VCCH m2_23680_n288167# sky130_fd_pr__cap_mim_m3_2_HYMU45
XXC4 m4_25183_n288425# VSS sky130_fd_pr__cap_mim_m3_2_4PHTN9
XXC5 VCCH m1_22999_n287228# sky130_fd_pr__cap_mim_m3_2_RQPX7Z
Xsky130_fd_pr__cap_mim_m3_2_4PHTN9_0 m2_24504_n284758# VSS sky130_fd_pr__cap_mim_m3_2_4PHTN9
Xsky130_fd_pr__cap_mim_m3_1_EEU5EF_0 VSS VT2 VT2 VSS sky130_fd_pr__cap_mim_m3_1_EEU5EF
XXC9 m2_24748_n284671# VSS sky130_fd_pr__cap_mim_m3_2_4PHTN9
Xsky130_fd_pr__cap_mim_m3_1_EEU5EF_1 VSS VT3 VT3 VSS sky130_fd_pr__cap_mim_m3_1_EEU5EF
Xsky130_fd_pr__cap_mim_m3_1_RRZ644_0 VCCH m2_23680_n288167# sky130_fd_pr__cap_mim_m3_1_RRZ644
XXM40 Td_Sd VCCL Td_Sd Td_Sd VCCL m2_24748_n284671# VCCL Td_Sd m2_24748_n284671# sky130_fd_pr__pfet_01v8_X6XW7S
XXM30 Td_L VSS VSS VSS m2_31884_n287663# sky130_fd_pr__nfet_01v8_5QNSAB
XXM31 VCCL Td_L VCCL VCCL Td_L m2_31884_n287663# VCCL VCCL m2_31884_n287663# sky130_fd_pr__pfet_01v8_X6XW7S
XXM20 vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__res_xhigh_po_0p69_KA8C77_2 m1_19785_n286949# m1_17211_n289349# m1_17679_n289349#
+ m1_22125_n286949# m1_20487_n289349# m1_16743_n289349# m1_19551_n289349# m1_18849_n286949#
+ m1_18381_n286949# m1_19551_n289349# m1_18849_n286949# m1_19083_n289349# m1_20019_n289349#
+ m1_16739_n286950# m1_21189_n286949# m1_20721_n286949# m1_16977_n286949# m1_20721_n286949#
+ m1_17211_n289349# m1_18147_n289349# m1_21891_n289349# m1_20955_n289349# m1_17679_n289349#
+ m1_16743_n289349# m1_17913_n286949# m1_18615_n289349# VSS m1_20019_n289349# m1_18381_n286949#
+ m1_17913_n286949# m1_19785_n286949# m1_21657_n286949# m1_21657_n286949# m1_21189_n286949#
+ m1_19317_n286949# m1_18147_n289349# m1_21423_n289349# m1_19083_n289349# m1_19317_n286949#
+ m1_20955_n289349# m1_21891_n289349# m1_21423_n289349# m1_20487_n289349# m1_18615_n289349#
+ m1_16977_n286949# m1_20253_n286949# m1_17445_n286949# m1_20253_n286949# m1_17445_n286949#
+ sky130_fd_pr__res_xhigh_po_0p69_KA8C77
XXM32 VSS VSS Td_S m4_25183_n288425# sky130_fd_pr__nfet_01v8_L9ESAD
XXM21 VSS m2_29342_n288187# VSS vbn1 vbn1 vbn1 vbn1 m2_29342_n288187# VSS m2_29342_n288187#
+ sky130_fd_pr__nfet_g5v0d10v5_XSEQJ6
XXM10 VT2 m2_29759_n286901# m2_30306_n287752# VCCL m2_30306_n287752# m2_29759_n286901#
+ sky130_fd_pr__pfet_01v8_6QC8WZ
XdelayPulse_digital_0 Td_Lb Td_Sd porbPre porPre Td_Sd Td_L VCCL VSS delayPulse_digital
Xsky130_fd_pr__res_xhigh_po_0p69_KA8C77_3 m1_20018_n283415# m1_16975_n285816# m1_17911_n285816#
+ m1_21890_n283415# m1_20719_n285816# m1_16739_n286950# m1_19783_n285816# m1_18614_n283415#
+ m1_18614_n283415# m1_19315_n285816# m1_19082_n283415# m1_18847_n285816# m1_20251_n285816#
+ m1_16742_n283415# m1_20954_n283415# m1_20954_n283415# m1_16742_n283415# m1_20486_n283415#
+ m1_17443_n285816# m1_17911_n285816# m1_21655_n285816# m1_21187_n285816# m1_17443_n285816#
+ m1_16975_n285816# m1_17678_n283415# m1_18379_n285816# VSS m1_19783_n285816# m1_18146_n283415#
+ m1_18146_n283415# m1_19550_n283415# m1_21890_n283415# m1_21422_n283415# m1_21422_n283415#
+ m1_19550_n283415# m1_18379_n285816# m1_21655_n285816# m1_19315_n285816# m1_19082_n283415#
+ m1_20719_n285816# VSS m1_21187_n285816# m1_20251_n285816# m1_18847_n285816# m1_17210_n283415#
+ m1_20486_n283415# m1_17678_n283415# m1_20018_n283415# m1_17210_n283415# sky130_fd_pr__res_xhigh_po_0p69_KA8C77
XXM33 VCCL Td_S VCCL VCCL m4_25183_n288425# Td_S m4_25183_n288425# sky130_fd_pr__pfet_01v8_U6B66J
XXM22[0] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[1] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[2] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[3] vbp2 vbp1 vbp2 vbp2 vbp1 VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM11 m2_23680_n288167# m2_24152_n287606# VCCH vbn1 sky130_fd_pr__pfet_g5v0d10v5_PQJ659
Xpor_output_buffer_0 VCCL porb VSS porbPre por_output_buffer
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_NZA8SD a_n699_n1416# a_n1529_984# a_n1861_n1416#
+ a_1293_n1416# a_463_n1416# a_1625_n1416# a_1293_984# a_297_984# a_n1861_984# a_n2157_n1546#
+ a_n865_984# a_n1363_n1416# a_n533_n1416# a_1127_n1416# a_1127_984# a_131_984# a_n35_n1416#
+ a_n1197_984# a_795_n1416# a_1957_n1416# a_1459_984# a_463_984# a_n1031_984# a_n1695_n1416#
+ a_297_n1416# a_n865_n1416# a_n2027_984# a_1459_n1416# a_629_n1416# a_1791_984# a_n35_984#
+ a_795_984# a_n1197_n1416# a_n367_984# a_n1363_984# a_n1529_n1416# a_n367_n1416#
+ a_1625_984# a_131_n1416# a_n2027_n1416# a_629_984# a_n201_984# a_n699_984# a_n1031_n1416#
+ a_n1695_984# a_1791_n1416# a_961_n1416# a_n201_n1416# a_1957_984# a_961_984# a_n533_984#
X0 a_131_984# a_131_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_1293_984# a_1293_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_n1031_984# a_n1031_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_629_984# a_629_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n1529_984# a_n1529_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_n699_984# a_n699_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_961_984# a_961_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_1459_984# a_1459_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n1861_984# a_n1861_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_n35_984# a_n35_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_n367_984# a_n367_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_1791_984# a_1791_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_1127_984# a_1127_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_297_984# a_297_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_n1197_984# a_n1197_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_1957_984# a_1957_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_n865_984# a_n865_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_1625_984# a_1625_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X18 a_n2027_984# a_n2027_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X19 a_n533_984# a_n533_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X20 a_795_984# a_795_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X21 a_n1695_984# a_n1695_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X22 a_n201_984# a_n201_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X23 a_463_984# a_463_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X24 a_n1363_984# a_n1363_n1416# a_n2157_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_D2SRCG a_n165_n1446# a_n35_n1316# a_n35_884#
X0 a_n35_884# a_n35_n1316# a_n165_n1446# sky130_fd_pr__res_xhigh_po_0p35 l=9
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_SZAJAG a_n699_n1416# a_463_n1416# a_297_984#
+ a_n865_984# a_n533_n1416# a_1127_n1416# a_1127_984# a_131_984# a_n35_n1416# a_n1197_984#
+ a_795_n1416# a_463_984# a_n1031_984# a_297_n1416# a_n865_n1416# a_629_n1416# a_n35_984#
+ a_795_984# a_n1197_n1416# a_n367_984# a_n367_n1416# a_n1327_n1546# a_131_n1416#
+ a_629_984# a_n201_984# a_n699_984# a_n1031_n1416# a_961_n1416# a_n201_n1416# a_961_984#
+ a_n533_984#
X0 a_131_984# a_131_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n1031_984# a_n1031_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_629_984# a_629_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n699_984# a_n699_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_961_984# a_961_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_n35_984# a_n35_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_n367_984# a_n367_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_1127_984# a_1127_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_297_984# a_297_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_n1197_984# a_n1197_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_n865_984# a_n865_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n533_984# a_n533_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_795_984# a_795_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_n201_984# a_n201_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_463_984# a_463_n1416# a_n1327_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_CZFQWY a_90_n309# a_n90_21# a_n148_n309# a_n282_n531#
+ a_n148_109# a_90_109# a_n90_n397#
X0 a_90_109# a_n90_21# a_n148_109# a_n282_n531# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
X1 a_90_n309# a_n90_n397# a_n148_n309# a_n282_n531# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
.ends

.subckt sky130_sw_ip__bgrref_por vbg por avdd dvdd porb porb_h[0] porb_h[1] avss dvss
Xx1 x1/Vinn x1/Vinp x2/din avdd dvdd avss comparator_final
Xx2 x2/din por vbg porb porb_h[0] porb_h[1] avdd dvdd dvss delayPulse_final
XXR1 m1_10262_n288829# m1_11092_n286429# m1_11258_n288829# m1_8270_n288829# m1_8934_n288829#
+ m1_7938_n288829# m1_8104_n286429# m1_9100_n286429# m1_11424_n286429# avss m1_10428_n286429#
+ m1_10926_n288829# m1_9930_n288829# m1_8270_n288829# m1_8436_n286429# m1_9432_n286429#
+ m1_9598_n288829# m1_10760_n286429# m1_8602_n288829# m1_7606_n288829# m1_8104_n286429#
+ m1_9100_n286429# m1_10428_n286429# m1_11258_n288829# m1_9266_n288829# m1_10262_n288829#
+ m1_11424_n286429# m1_7938_n288829# m1_8934_n288829# m1_7772_n286429# m1_9432_n286429#
+ m1_8768_n286429# m1_10594_n288829# m1_9764_n286429# m1_10760_n286429# m1_10926_n288829#
+ m1_9930_n288829# m1_7772_n286429# m1_9266_n288829# x1/Vinn m1_8768_n286429# m1_9764_n286429#
+ m1_10096_n286429# m1_10594_n288829# m1_11092_n286429# m1_7606_n288829# m1_8602_n288829#
+ m1_9598_n288829# avss m1_8436_n286429# m1_10096_n286429# sky130_fd_pr__res_xhigh_po_0p35_NZA8SD
XXR10 avss x1/Vinn x1/Vinp sky130_fd_pr__res_xhigh_po_0p35_D2SRCG
XXR12 m1_14304_n288829# m1_13302_n288829# m1_13468_n286429# m1_14470_n286429# m1_14304_n288829#
+ m1_12634_n288829# x1/Vinp m1_13468_n286429# m1_13636_n288829# m1_14804_n286429#
+ m1_12968_n288829# m1_13134_n286429# m1_14804_n286429# m1_13302_n288829# m1_14638_n288829#
+ m1_12968_n288829# m1_13802_n286429# m1_12800_n286429# m1_14983_n288829# m1_14136_n286429#
+ m1_13970_n288829# avss m1_13636_n288829# m1_13134_n286429# m1_13802_n286429# m1_14470_n286429#
+ m1_14638_n288829# m1_12634_n288829# m1_13970_n288829# m1_12800_n286429# m1_14136_n286429#
+ sky130_fd_pr__res_xhigh_po_0p35_SZAJAG
XXM2 avdd avdd m1_14983_n288829# avss m1_14983_n288829# avdd avdd sky130_fd_pr__nfet_05v0_nvt_CZFQWY
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9992MR__0 a_50_n136# a_n108_n136# a_n50_n162#
+ w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt poly_res_200ohm a_n414_974# a_n414_n76#
X0 a_n414_974# a_n414_n76# sky130_fd_pr__res_generic_po w=0.71 l=2.96
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0 a_n108_n34# a_n50_n122# a_50_n34# VSUBS
X0 a_50_n34# a_n50_n122# a_n108_n34# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.1885 pd=1.88 as=0.1885 ps=1.88 w=0.65 l=0.5
.ends

.subckt rheo_3v_cell_top m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ w_318_892# m1_290_1114# poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125#
+ m4_97_801# m1_821_212# m4_97_1059# m1_814_483# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_1 m1_824_799# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt rheo_3v_cell m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_290_1114#
+ poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125# m1_821_212# m1_824_799#
+ m1_814_483# poly_res_200ohm_1/a_n414_974# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# w_316_892# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt rheo_3v_column rheo_3v_cell_top_0/m4_97_1059# b3b b0_uq14 b0_uq3 b2b_uq1 dum1_out
+ b0_uq2 rheo_3v_cell_0[1]/w_316_892# b0b_uq14 b3 rheo_3v_cell_top_0/m1_290_591# b1_uq6
+ b0b_uq9 rheo_3v_cell_0[5]/w_316_892# b0_uq13 b0b_uq12 b1 rheo_3v_cell_0[6]/w_316_892#
+ b0b_uq8 dum0_in b0b_uq7 b2 b1_uq3 b0_uq0 b0b_uq6 b1_uq2 rheo_3v_cell_top_0/m1_290_1114#
+ b1_uq1 b1_uq5 b1_uq0 b3_uq0 b3b_uq0 b1_uq4 b0b_uq5 rheo_3v_cell_0[4]/w_316_892#
+ b0_uq5 m2_801_196# rheo_3v_cell_0[7]/w_316_892# b0b_uq0 b0b_uq13 b0_uq4 b0b_uq4
+ out_5 b0_uq11 b2b_uq0 out_4 b4 b0_uq10 rheo_3v_cell_0[3]/w_316_892# b2_uq2 b0b_uq3
+ b2_uq1 b0_uq12 m2_801_13759# res0_in b0b_uq1 b0b_uq2 b1b_uq3 b1b_uq4 b1b_uq6 b1b_uq2
+ b4b b1b_uq1 b2b_uq2 b1b_uq0 b1b_uq5 m2_791_1314# b2_uq0 b0b_uq11 rheo_3v_cell_0[2]/w_316_892#
+ b0_uq9 b0b b0_uq1 res1_out b0_uq8 rheo_3v_cell_top_0/m4_97_801# b0_uq6 b0b_uq10
+ m2_791_14877# b1b b0_uq7 b0 b2b VSUBS
Xrheo_3v_cell_top_0 b0_uq14 rheo_3v_cell_0[7]/w_316_892# out_4 out_5 res1_in m2_801_13759#
+ rheo_3v_cell_top_0/m1_290_1114# VSUBS out0_0_3 out1_0_0 b0b_uq13 rheo_3v_cell_top_0/m4_97_801#
+ out1_1_0 rheo_3v_cell_top_0/m4_97_1059# b1_uq6 rheo_3v_cell_0[7]/m1_824_799# out1_0_0
+ rheo_3v_cell_top_0/m1_155_n223# b0b_uq14 b1b_uq6 rheo_3v_cell_top_0/m1_290_591#
+ b0_uq13 rheo_3v_cell_top
Xrheo_3v_cell_0[0] m2_791_1314# m2_801_196# m2_328_1119# m2_328_1119# m2_791_1314#
+ VSUBS m2_449_485# m2_328_1119# m2_801_196# m2_449_485# res1_out VSUBS res0_in dum1_out
+ m2_449_485# dum0_in VSUBS m2_791_1314# m2_801_196# VSUBS VSUBS rheo_3v_cell
Xrheo_3v_cell_0[1] b0b m2_791_1314# out0_0_0 out0_1_0 b1b_uq0 VSUBS out0_0_0 out1_0_3
+ b0_uq0 out_3 rheo_3v_cell_0[1]/m1_824_799# b4b rheo_3v_cell_0[2]/m1_155_n223# res1_out
+ out_4 res0_in b0 rheo_3v_cell_0[1]/w_316_892# b4 b1_uq0 b0b_uq0 rheo_3v_cell
Xrheo_3v_cell_0[2] b0_uq2 rheo_3v_cell_0[1]/w_316_892# out0_2 out0_1_0 b2b_uq0 VSUBS
+ out0_0_0 out1_0_3 b0b_uq1 out1_1_1 rheo_3v_cell_0[2]/m1_824_799# b1b rheo_3v_cell_0[3]/m1_155_n223#
+ rheo_3v_cell_0[1]/m1_824_799# out1_0_3 rheo_3v_cell_0[2]/m1_155_n223# b0b_uq2 rheo_3v_cell_0[2]/w_316_892#
+ b1 b2_uq0 b0_uq1 rheo_3v_cell
Xrheo_3v_cell_0[3] b0b_uq4 rheo_3v_cell_0[2]/w_316_892# out0_0_1 out0_1_0 b1_uq1 VSUBS
+ out0_0_1 out1_0_2 b0_uq3 out1_1_1 rheo_3v_cell_0[3]/m1_824_799# b2b rheo_3v_cell_0[4]/m1_155_n223#
+ rheo_3v_cell_0[2]/m1_824_799# out1_2 rheo_3v_cell_0[3]/m1_155_n223# b0_uq4 rheo_3v_cell_0[3]/w_316_892#
+ b2 b1b_uq1 b0b_uq3 rheo_3v_cell
Xrheo_3v_cell_0[4] b0_uq6 rheo_3v_cell_0[3]/w_316_892# out_3 out0_2 b3b_uq0 VSUBS
+ out0_0_1 out1_0_2 b0b_uq5 out1_1_1 rheo_3v_cell_0[4]/m1_824_799# b1_uq2 rheo_3v_cell_0[5]/m1_155_n223#
+ rheo_3v_cell_0[3]/m1_824_799# out1_0_2 rheo_3v_cell_0[4]/m1_155_n223# b0b_uq6 rheo_3v_cell_0[4]/w_316_892#
+ b1b_uq2 b3_uq0 b0_uq5 rheo_3v_cell
Xrheo_3v_cell_0[5] b0b_uq8 rheo_3v_cell_0[4]/w_316_892# out0_0_2 out0_1_1 b1b_uq3
+ VSUBS out0_0_2 out1_0_1 b0_uq7 out1_2 rheo_3v_cell_0[5]/m1_824_799# b3b rheo_3v_cell_0[6]/m1_155_n223#
+ rheo_3v_cell_0[4]/m1_824_799# out_3 rheo_3v_cell_0[5]/m1_155_n223# b0_uq8 rheo_3v_cell_0[5]/w_316_892#
+ b3 b1_uq3 b0b_uq7 rheo_3v_cell
Xrheo_3v_cell_0[6] b0_uq10 rheo_3v_cell_0[5]/w_316_892# out0_2 out0_1_1 b2_uq1 VSUBS
+ out0_0_2 out1_0_1 b0b_uq9 out1_1_0 rheo_3v_cell_0[6]/m1_824_799# b1b_uq4 rheo_3v_cell_0[7]/m1_155_n223#
+ rheo_3v_cell_0[5]/m1_824_799# out1_0_1 rheo_3v_cell_0[6]/m1_155_n223# b0b_uq10 rheo_3v_cell_0[6]/w_316_892#
+ b1_uq4 b2b_uq1 b0_uq9 rheo_3v_cell
Xrheo_3v_cell_0[7] b0b_uq12 rheo_3v_cell_0[6]/w_316_892# out0_0_3 out0_1_1 b1_uq5
+ VSUBS out0_0_3 out1_0_0 b0_uq11 out1_1_0 rheo_3v_cell_0[7]/m1_824_799# b2_uq2 rheo_3v_cell_top_0/m1_155_n223#
+ rheo_3v_cell_0[6]/m1_824_799# out1_2 rheo_3v_cell_0[7]/m1_155_n223# b0_uq12 rheo_3v_cell_0[7]/w_316_892#
+ b2b_uq2 b1b_uq5 b0b_uq11 rheo_3v_cell
Xrheo_3v_cell_1 m2_791_14877# m2_801_13759# m2_330_14682# m2_330_14682# m2_791_14877#
+ VSUBS m2_449_14048# m2_330_14682# m2_801_13759# m2_449_14048# dum0_out VSUBS dum0_out
+ res1_in m2_449_14048# res1_in VSUBS m2_791_14877# m2_801_13759# VSUBS VSUBS rheo_3v_cell
.ends

.subckt rheo_3v_cell_odd m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_290_1114#
+ poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125# m1_821_212# m1_824_799#
+ m1_814_483# poly_res_200ohm_1/a_n414_974# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# w_316_892# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt rheo_3v_column_odd rheo_3v_cell_top_0/m4_97_1059# m3_31_13582# res_in0 b0_uq14
+ b2b_uq2 b0_uq12 b0_uq6 rheo_3v_cell_0[1]/w_316_892# b0b_uq14 b1_uq6 rheo_3v_cell_0[0]/w_316_892#
+ b0_uq1 b0_uq13 b0b_uq12 b1 in_5 b0b_uq11 b3 b0b_uq10 b0_uq3 b3b b1_uq1 m3_30_13212#
+ b0_uq2 b0b_uq3 b2b_uq1 b0_uq0 b0b_uq9 rheo_3v_cell_0[4]/w_316_892# b0b_uq2 rheo_3v_cell_odd_0/w_316_892#
+ rheo_3v_cell_0[5]/w_316_892# b0b_uq1 b0b_uq13 b0b_uq8 b3b_uq0 b1_uq2 b4 b2 out_5
+ b1_uq3 dum_in0 res_out1 rheo_3v_cell_0[3]/w_316_892# b2_uq2 b0b_uq7 b1_uq5 b4b out4
+ b1b_uq5 b2_uq1 b1_uq4 m2_801_196# m2_791_14877# m2_801_13759# b1b_uq4 b0b_uq6 b0b_uq5
+ b0 b2_uq0 b1b_uq3 b1b_uq6 b1b_uq2 b0b_uq4 b1b_uq1 b1b_uq0 b0_uq11 b2b_uq0 b3_uq0
+ b1_uq0 rheo_3v_cell_0[2]/w_316_892# b0_uq9 dum_out1 b0_uq5 b0b b0b_uq0 b0_uq8 rheo_3v_cell_top_0/m4_97_801#
+ b0_uq10 m2_791_1314# b1b VSUBS b0_uq7 b0_uq4 b2b
Xrheo_3v_cell_2 m2_791_14877# m2_801_13759# m2_331_14682# m2_331_14682# m2_791_14877#
+ VSUBS m2_458_14048# m2_331_14682# m2_801_13759# m2_458_14048# dum_out0 VSUBS dum_out0
+ res_in1 m2_458_14048# res_in1 VSUBS m2_791_14877# m2_801_13759# VSUBS VSUBS rheo_3v_cell
Xrheo_3v_cell_odd_0 b0b m2_791_1314# out0_0_0 out0_1_0 b1b_uq0 VSUBS out0_0_0 out1_0_3
+ b0_uq0 out_3 rheo_3v_cell_odd_0/m1_824_799# b4 rheo_3v_cell_0[0]/m1_155_n223# res_out1
+ out4 res_in0 b0 rheo_3v_cell_odd_0/w_316_892# b4b b1_uq0 b0b_uq0 rheo_3v_cell_odd
Xrheo_3v_cell_top_0 b0_uq14 rheo_3v_cell_0[5]/w_316_892# in_5 out_5 res_in1 m2_801_13759#
+ m3_31_13582# VSUBS out0_0_3 out1_0_0 b0b_uq13 rheo_3v_cell_top_0/m4_97_801# out1_1_0
+ rheo_3v_cell_top_0/m4_97_1059# b1_uq6 rheo_3v_cell_0[5]/m1_824_799# out1_0_0 rheo_3v_cell_top_0/m1_155_n223#
+ b0b_uq14 b1b_uq6 m3_30_13212# b0_uq13 rheo_3v_cell_top
Xrheo_3v_cell_0[0] b0_uq2 rheo_3v_cell_odd_0/w_316_892# out0_2 out0_1_0 b2b_uq0 VSUBS
+ out0_0_0 out1_0_3 b0b_uq1 out1_1_1 rheo_3v_cell_0[0]/m1_824_799# b1b rheo_3v_cell_0[1]/m1_155_n223#
+ rheo_3v_cell_odd_0/m1_824_799# out1_0_3 rheo_3v_cell_0[0]/m1_155_n223# b0b_uq2 rheo_3v_cell_0[0]/w_316_892#
+ b1 b2_uq0 b0_uq1 rheo_3v_cell
Xrheo_3v_cell_0[1] b0b_uq4 rheo_3v_cell_0[0]/w_316_892# out0_0_1 out0_1_0 b1_uq1 VSUBS
+ out0_0_1 out1_0_2 b0_uq3 out1_1_1 rheo_3v_cell_0[1]/m1_824_799# b2b rheo_3v_cell_0[2]/m1_155_n223#
+ rheo_3v_cell_0[0]/m1_824_799# out1_2 rheo_3v_cell_0[1]/m1_155_n223# b0_uq4 rheo_3v_cell_0[1]/w_316_892#
+ b2 b1b_uq1 b0b_uq3 rheo_3v_cell
Xrheo_3v_cell_0[2] b0_uq6 rheo_3v_cell_0[1]/w_316_892# out_3 out0_2 b3b_uq0 VSUBS
+ out0_0_1 out1_0_2 b0b_uq5 out1_1_1 rheo_3v_cell_0[2]/m1_824_799# b1_uq2 rheo_3v_cell_0[3]/m1_155_n223#
+ rheo_3v_cell_0[1]/m1_824_799# out1_0_2 rheo_3v_cell_0[2]/m1_155_n223# b0b_uq6 rheo_3v_cell_0[2]/w_316_892#
+ b1b_uq2 b3_uq0 b0_uq5 rheo_3v_cell
Xrheo_3v_cell_0[3] b0b_uq8 rheo_3v_cell_0[2]/w_316_892# out0_0_2 m3_296_8710# b1b_uq3
+ VSUBS out0_0_2 out1_0_1 b0_uq7 out1_2 rheo_3v_cell_0[3]/m1_824_799# b3b rheo_3v_cell_0[4]/m1_155_n223#
+ rheo_3v_cell_0[2]/m1_824_799# out_3 rheo_3v_cell_0[3]/m1_155_n223# b0_uq8 rheo_3v_cell_0[3]/w_316_892#
+ b3 b1_uq3 b0b_uq7 rheo_3v_cell
Xrheo_3v_cell_0[4] b0_uq10 rheo_3v_cell_0[3]/w_316_892# out0_2 m3_296_8710# b2_uq1
+ VSUBS out0_0_2 out1_0_1 b0b_uq9 out1_1_0 rheo_3v_cell_0[4]/m1_824_799# b1b_uq4 rheo_3v_cell_0[5]/m1_155_n223#
+ rheo_3v_cell_0[3]/m1_824_799# out1_0_1 rheo_3v_cell_0[4]/m1_155_n223# b0b_uq10 rheo_3v_cell_0[4]/w_316_892#
+ b1_uq4 b2b_uq1 b0_uq9 rheo_3v_cell
Xrheo_3v_cell_0[5] b0b_uq12 rheo_3v_cell_0[4]/w_316_892# out0_0_3 m3_296_8710# b1_uq5
+ VSUBS out0_0_3 out1_0_0 b0_uq11 out1_1_0 rheo_3v_cell_0[5]/m1_824_799# b2_uq2 rheo_3v_cell_top_0/m1_155_n223#
+ rheo_3v_cell_0[4]/m1_824_799# out1_2 rheo_3v_cell_0[5]/m1_155_n223# b0_uq12 rheo_3v_cell_0[5]/w_316_892#
+ b2b_uq2 b1b_uq5 b0b_uq11 rheo_3v_cell
Xrheo_3v_cell_1 m2_791_1314# m2_801_196# m2_329_1119# m2_329_1119# m2_791_1314# VSUBS
+ m2_457_485# m2_329_1119# m2_801_196# m2_457_485# res_out1 VSUBS res_in0 dum_out1
+ m2_457_485# dum_in0 VSUBS m2_791_1314# m2_801_196# VSUBS VSUBS rheo_3v_cell
.ends

.subckt rheo_3v_cell_dummy m4_99_18# w_318_n275# m4_99_276# m4_99_801# poly_res_200ohm_1/VSUBS
+ m4_99_930# m1_824_799# poly_res_200ohm_1/a_n414_974# m4_99_405# m4_99_1059# poly_res_200ohm_0/a_n414_n76#
+ m4_99_672# m1_155_n223# w_316_892# m4_99_147#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_387_847# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_545_212# m1_545_212# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# poly_res_200ohm_1/VSUBS m1_387_847#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_387_847# poly_res_200ohm_1/VSUBS m1_824_799#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# poly_res_200ohm_1/VSUBS m1_545_212#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_545_212# poly_res_200ohm_1/VSUBS m1_545_212#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt rheo_3v_column_dummy rheo_3v_cell_dummy_0[7]/m4_99_930# rheo_3v_cell_dummy_0[7]/m4_99_1059#
+ rheo_3v_cell_dummy_0[2]/m4_99_1059# rheo_3v_cell_dummy_0[8]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_930#
+ rheo_3v_cell_dummy_0[0]/m4_99_405# rheo_3v_cell_dummy_0[9]/m4_99_930# rheo_3v_cell_dummy_0[1]/m4_99_405#
+ rheo_3v_cell_dummy_0[2]/m4_99_405# rheo_3v_cell_dummy_0[0]/m4_99_672# rheo_3v_cell_dummy_0[9]/m4_99_18#
+ rheo_3v_cell_dummy_0[1]/m4_99_672# rheo_3v_cell_dummy_0[3]/m4_99_405# rheo_3v_cell_dummy_0[2]/m4_99_672#
+ rheo_3v_cell_dummy_0[4]/m4_99_405# rheo_3v_cell_dummy_0[5]/m4_99_405# rheo_3v_cell_dummy_0[3]/m4_99_672#
+ rheo_3v_cell_dummy_0[6]/m4_99_405# rheo_3v_cell_dummy_0[4]/m4_99_672# rheo_3v_cell_dummy_0[3]/w_316_892#
+ rheo_3v_cell_dummy_0[5]/m4_99_672# rheo_3v_cell_dummy_0[7]/m4_99_405# rheo_3v_cell_dummy_0[6]/m4_99_1059#
+ rheo_3v_cell_dummy_0[1]/m4_99_1059# rheo_3v_cell_dummy_0[8]/m4_99_405# rheo_3v_cell_dummy_0[6]/m4_99_672#
+ rheo_3v_cell_dummy_0[7]/m4_99_672# rheo_3v_cell_dummy_0[9]/m4_99_405# rheo_3v_cell_dummy_0[2]/w_316_892#
+ rheo_3v_cell_dummy_0[8]/m4_99_672# rheo_3v_cell_dummy_0[0]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_147#
+ rheo_3v_cell_dummy_0[7]/w_316_892# rheo_3v_cell_dummy_0[9]/m4_99_672# rheo_3v_cell_dummy_0[8]/w_316_892#
+ rheo_3v_cell_dummy_0[1]/m4_99_147# rheo_3v_cell_dummy_0[9]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_147#
+ rheo_3v_cell_dummy_0[3]/m4_99_147# rheo_3v_cell_dummy_0[1]/m4_99_18# rheo_3v_cell_dummy_0[4]/m4_99_147#
+ rheo_3v_cell_dummy_0[5]/m4_99_147# rheo_3v_cell_dummy_0[5]/m4_99_1059# rheo_3v_cell_dummy_0[0]/m4_99_1059#
+ rheo_3v_cell_dummy_0[6]/m4_99_147# rheo_3v_cell_dummy_0[6]/w_316_892# rheo_3v_cell_dummy_0[7]/m4_99_147#
+ rheo_3v_cell_dummy_0[1]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_147#
+ rheo_3v_cell_dummy_0[9]/m4_99_147# rheo_3v_cell_dummy_0[3]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_276#
+ rheo_3v_cell_dummy_0[0]/m4_99_801# rheo_3v_cell_dummy_0[1]/m4_99_276# rheo_3v_cell_dummy_0[9]/m4_99_1059#
+ rheo_3v_cell_dummy_0[1]/m4_99_801# rheo_3v_cell_dummy_0[4]/m4_99_1059# rheo_3v_cell_dummy_0[2]/m4_99_276#
+ rheo_3v_cell_dummy_0[2]/m4_99_801# rheo_3v_cell_dummy_0[3]/m4_99_276# rheo_3v_cell_dummy_0[3]/m4_99_801#
+ rheo_3v_cell_dummy_0[5]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_18# rheo_3v_cell_dummy_0[4]/m4_99_276#
+ rheo_3v_cell_dummy_0[0]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_801# rheo_3v_cell_dummy_0[5]/m4_99_276#
+ rheo_3v_cell_dummy_0[5]/m4_99_801# rheo_3v_cell_dummy_0[6]/m4_99_276# rheo_3v_cell_dummy_0[6]/m4_99_801#
+ rheo_3v_cell_dummy_0[7]/m4_99_276# rheo_3v_cell_dummy_0[7]/m4_99_801# rheo_3v_cell_dummy_0[8]/m4_99_276#
+ rheo_3v_cell_dummy_0[5]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_801# rheo_3v_cell_dummy_0[9]/m4_99_276#
+ rheo_3v_cell_dummy_0[9]/m4_99_801# rheo_3v_cell_dummy_0[8]/m4_99_1059# rheo_3v_cell_dummy_0[3]/m4_99_1059#
+ rheo_3v_cell_dummy_0[6]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_930# rheo_3v_cell_dummy_0[4]/w_316_892#
+ rheo_3v_cell_dummy_0[0]/w_318_n275# rheo_3v_cell_dummy_0[1]/m4_99_930# rheo_3v_cell_dummy_0[2]/m4_99_930#
+ m1_988_1608# rheo_3v_cell_dummy_0[3]/m4_99_930# rheo_3v_cell_dummy_0[7]/m4_99_18#
+ m1_n18_1607# rheo_3v_cell_dummy_0[4]/m4_99_930# m1_938_45# rheo_3v_cell_dummy_0[5]/m4_99_930#
+ rheo_3v_cell_dummy_0[6]/m4_99_930# m1_n18_45# VSUBS
Xrheo_3v_cell_dummy_0[0] rheo_3v_cell_dummy_0[0]/m4_99_18# rheo_3v_cell_dummy_0[0]/w_318_n275#
+ rheo_3v_cell_dummy_0[0]/m4_99_276# rheo_3v_cell_dummy_0[0]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[0]/m4_99_930#
+ m1_988_1608# m1_n18_1607# rheo_3v_cell_dummy_0[0]/m4_99_405# rheo_3v_cell_dummy_0[0]/m4_99_1059#
+ m1_938_45# rheo_3v_cell_dummy_0[0]/m4_99_672# m1_n18_45# rheo_3v_cell_dummy_0[0]/w_316_892#
+ rheo_3v_cell_dummy_0[0]/m4_99_147# rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[1] rheo_3v_cell_dummy_0[1]/m4_99_18# rheo_3v_cell_dummy_0[0]/w_316_892#
+ rheo_3v_cell_dummy_0[1]/m4_99_276# rheo_3v_cell_dummy_0[1]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[1]/m4_99_930#
+ rheo_3v_cell_dummy_0[1]/m1_824_799# rheo_3v_cell_dummy_0[2]/m1_155_n223# rheo_3v_cell_dummy_0[1]/m4_99_405#
+ rheo_3v_cell_dummy_0[1]/m4_99_1059# m1_988_1608# rheo_3v_cell_dummy_0[1]/m4_99_672#
+ m1_n18_1607# rheo_3v_cell_dummy_0[1]/w_316_892# rheo_3v_cell_dummy_0[1]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[2] rheo_3v_cell_dummy_0[2]/m4_99_18# rheo_3v_cell_dummy_0[1]/w_316_892#
+ rheo_3v_cell_dummy_0[2]/m4_99_276# rheo_3v_cell_dummy_0[2]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[2]/m4_99_930#
+ rheo_3v_cell_dummy_0[2]/m1_824_799# rheo_3v_cell_dummy_0[3]/m1_155_n223# rheo_3v_cell_dummy_0[2]/m4_99_405#
+ rheo_3v_cell_dummy_0[2]/m4_99_1059# rheo_3v_cell_dummy_0[1]/m1_824_799# rheo_3v_cell_dummy_0[2]/m4_99_672#
+ rheo_3v_cell_dummy_0[2]/m1_155_n223# rheo_3v_cell_dummy_0[2]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[3] rheo_3v_cell_dummy_0[3]/m4_99_18# rheo_3v_cell_dummy_0[2]/w_316_892#
+ rheo_3v_cell_dummy_0[3]/m4_99_276# rheo_3v_cell_dummy_0[3]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[3]/m4_99_930#
+ rheo_3v_cell_dummy_0[3]/m1_824_799# rheo_3v_cell_dummy_0[4]/m1_155_n223# rheo_3v_cell_dummy_0[3]/m4_99_405#
+ rheo_3v_cell_dummy_0[3]/m4_99_1059# rheo_3v_cell_dummy_0[2]/m1_824_799# rheo_3v_cell_dummy_0[3]/m4_99_672#
+ rheo_3v_cell_dummy_0[3]/m1_155_n223# rheo_3v_cell_dummy_0[3]/w_316_892# rheo_3v_cell_dummy_0[3]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[4] rheo_3v_cell_dummy_0[4]/m4_99_18# rheo_3v_cell_dummy_0[3]/w_316_892#
+ rheo_3v_cell_dummy_0[4]/m4_99_276# rheo_3v_cell_dummy_0[4]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[4]/m4_99_930#
+ rheo_3v_cell_dummy_0[4]/m1_824_799# rheo_3v_cell_dummy_0[5]/m1_155_n223# rheo_3v_cell_dummy_0[4]/m4_99_405#
+ rheo_3v_cell_dummy_0[4]/m4_99_1059# rheo_3v_cell_dummy_0[3]/m1_824_799# rheo_3v_cell_dummy_0[4]/m4_99_672#
+ rheo_3v_cell_dummy_0[4]/m1_155_n223# rheo_3v_cell_dummy_0[4]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[5] rheo_3v_cell_dummy_0[5]/m4_99_18# rheo_3v_cell_dummy_0[4]/w_316_892#
+ rheo_3v_cell_dummy_0[5]/m4_99_276# rheo_3v_cell_dummy_0[5]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[5]/m4_99_930#
+ rheo_3v_cell_dummy_0[5]/m1_824_799# rheo_3v_cell_dummy_0[6]/m1_155_n223# rheo_3v_cell_dummy_0[5]/m4_99_405#
+ rheo_3v_cell_dummy_0[5]/m4_99_1059# rheo_3v_cell_dummy_0[4]/m1_824_799# rheo_3v_cell_dummy_0[5]/m4_99_672#
+ rheo_3v_cell_dummy_0[5]/m1_155_n223# rheo_3v_cell_dummy_0[5]/w_316_892# rheo_3v_cell_dummy_0[5]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[6] rheo_3v_cell_dummy_0[6]/m4_99_18# rheo_3v_cell_dummy_0[5]/w_316_892#
+ rheo_3v_cell_dummy_0[6]/m4_99_276# rheo_3v_cell_dummy_0[6]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[6]/m4_99_930#
+ rheo_3v_cell_dummy_0[6]/m1_824_799# rheo_3v_cell_dummy_0[7]/m1_155_n223# rheo_3v_cell_dummy_0[6]/m4_99_405#
+ rheo_3v_cell_dummy_0[6]/m4_99_1059# rheo_3v_cell_dummy_0[5]/m1_824_799# rheo_3v_cell_dummy_0[6]/m4_99_672#
+ rheo_3v_cell_dummy_0[6]/m1_155_n223# rheo_3v_cell_dummy_0[6]/w_316_892# rheo_3v_cell_dummy_0[6]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[7] rheo_3v_cell_dummy_0[7]/m4_99_18# rheo_3v_cell_dummy_0[6]/w_316_892#
+ rheo_3v_cell_dummy_0[7]/m4_99_276# rheo_3v_cell_dummy_0[7]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[7]/m4_99_930#
+ rheo_3v_cell_dummy_0[7]/m1_824_799# rheo_3v_cell_dummy_0[8]/m1_155_n223# rheo_3v_cell_dummy_0[7]/m4_99_405#
+ rheo_3v_cell_dummy_0[7]/m4_99_1059# rheo_3v_cell_dummy_0[6]/m1_824_799# rheo_3v_cell_dummy_0[7]/m4_99_672#
+ rheo_3v_cell_dummy_0[7]/m1_155_n223# rheo_3v_cell_dummy_0[7]/w_316_892# rheo_3v_cell_dummy_0[7]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[8] rheo_3v_cell_dummy_0[8]/m4_99_18# rheo_3v_cell_dummy_0[7]/w_316_892#
+ rheo_3v_cell_dummy_0[8]/m4_99_276# rheo_3v_cell_dummy_0[8]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[8]/m4_99_930#
+ m1_36_13186# m1_36_13186# rheo_3v_cell_dummy_0[8]/m4_99_405# rheo_3v_cell_dummy_0[8]/m4_99_1059#
+ rheo_3v_cell_dummy_0[7]/m1_824_799# rheo_3v_cell_dummy_0[8]/m4_99_672# rheo_3v_cell_dummy_0[8]/m1_155_n223#
+ rheo_3v_cell_dummy_0[8]/w_316_892# rheo_3v_cell_dummy_0[8]/m4_99_147# rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[9] rheo_3v_cell_dummy_0[9]/m4_99_18# rheo_3v_cell_dummy_0[8]/w_316_892#
+ rheo_3v_cell_dummy_0[9]/m4_99_276# rheo_3v_cell_dummy_0[9]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[9]/m4_99_930#
+ m1_28_15111# m1_28_15111# rheo_3v_cell_dummy_0[9]/m4_99_405# rheo_3v_cell_dummy_0[9]/m4_99_1059#
+ m1_36_13186# rheo_3v_cell_dummy_0[9]/m4_99_672# m1_36_13186# rheo_3v_cell_dummy_0[9]/w_316_892#
+ rheo_3v_cell_dummy_0[9]/m4_99_147# rheo_3v_cell_dummy
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.20625 pd=2.05 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.1575 ps=1.17 w=0.75 l=0.5
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_4AXGXB__0 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt rheo_level_shifter dvdd avdd bitb_out bit_out bit_in agnd
Xsky130_fd_sc_hvl__inv_8_1 bitb_out agnd agnd avdd avdd bit_out sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 bit_in dvdd agnd avdd avdd sky130_fd_sc_hvl__inv_2_0/A
+ avdd agnd agnd sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_4AXGXB_0 agnd bit_in sky130_fd_pr__diode_pw2nd_05v5_4AXGXB__0
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A agnd agnd avdd avdd bitb_out
+ sky130_fd_sc_hvl__inv_8
.ends

.subckt rheo_level_shifter_array rheo_level_shifter_0[0]/bit_in rheo_level_shifter_0[3]/bit_out
+ rheo_level_shifter_0[3]/bitb_out rheo_level_shifter_0[4]/bit_in rheo_level_shifter_0[0]/bit_out
+ rheo_level_shifter_0[4]/bitb_out rheo_level_shifter_0[7]/bit_out rheo_level_shifter_0[1]/bit_in
+ rheo_level_shifter_0[0]/bitb_out rheo_level_shifter_0[5]/bit_in rheo_level_shifter_0[4]/bit_out
+ rheo_level_shifter_0[7]/bitb_out rheo_level_shifter_0[1]/bit_out rheo_level_shifter_0[5]/bitb_out
+ rheo_level_shifter_0[1]/bitb_out rheo_level_shifter_0[6]/bit_in rheo_level_shifter_0[2]/bit_in
+ rheo_level_shifter_0[5]/bit_out rheo_level_shifter_0[6]/bitb_out rheo_level_shifter_0[2]/bit_out
+ rheo_level_shifter_0[2]/bitb_out rheo_level_shifter_0[3]/bit_in rheo_level_shifter_0[7]/bit_in
+ rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd rheo_level_shifter_0[6]/bit_out
+ VSUBS
Xrheo_level_shifter_0[0] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[0]/bitb_out rheo_level_shifter_0[0]/bit_out rheo_level_shifter_0[0]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[1] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[1]/bitb_out rheo_level_shifter_0[1]/bit_out rheo_level_shifter_0[1]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[2] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[2]/bitb_out rheo_level_shifter_0[2]/bit_out rheo_level_shifter_0[2]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[3] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[3]/bitb_out rheo_level_shifter_0[3]/bit_out rheo_level_shifter_0[3]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[4] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[4]/bitb_out rheo_level_shifter_0[4]/bit_out rheo_level_shifter_0[4]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[5] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[5]/bitb_out rheo_level_shifter_0[5]/bit_out rheo_level_shifter_0[5]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[6] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[6]/bitb_out rheo_level_shifter_0[6]/bit_out rheo_level_shifter_0[6]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[7] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[7]/bitb_out rheo_level_shifter_0[7]/bit_out rheo_level_shifter_0[7]/bit_in
+ VSUBS rheo_level_shifter
.ends

.subckt sky130_ef_ip__rheostat_8bit b0 b1 b2 b3 b4 b5 b6 b7 out vdd dvdd Vhigh Vlow
+ vss dvss
Xrheo_3v_column_0 b5a b3a b0b b0b b2a rheo_3v_column_0/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_0/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_1/out_5
+ b0b b2a rheo_3v_column_0/out_4 b4a b0b vdd b2b b0a b2b b0b vdd Vhigh b0a b0a b1a
+ b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_0/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_1 b5a b3a b0b b0b b2a rheo_3v_column_1/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_1/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_1/out_5
+ b0b b2a rheo_3v_column_1/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_1/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_1/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_2 b5a b3a b0b b0b b2a rheo_3v_column_2/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_2/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_3/out_5
+ b0b b2a rheo_3v_column_2/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_2/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_2/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_3 b5a b3a b0b b0b b2a rheo_3v_column_3/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_3/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_3/out_5
+ b0b b2a rheo_3v_column_3/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_3/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_3/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_4 b5a b3a b0b b0b b2a rheo_3v_column_4/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_4/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_5/out_5
+ b0b b2a rheo_3v_column_4/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_4/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_4/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_5 b5a b3a b0b b0b b2a rheo_3v_column_5/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_5/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_5/out_5
+ b0b b2a rheo_3v_column_5/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_5/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_5/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_6 b5a b3a b0b b0b b2a rheo_3v_column_6/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_6/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_7/out_5
+ b0b b2a rheo_3v_column_6/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_6/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_6/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_7 b5a b3a b0b b0b b2a rheo_3v_column_7/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_7/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_7/out_5
+ b0b b2a rheo_3v_column_7/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_7/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_7/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_odd_0 b5a b6b rheo_3v_column_0/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b6a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_1/out_5 b1b
+ rheo_3v_column_0/dum1_out rheo_3v_column_1/res0_in vdd b2b b0a b1b b4b rheo_3v_column_0/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_1/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_1 b5a b7b rheo_3v_column_1/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b7a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b out b1b rheo_3v_column_1/dum1_out
+ rheo_3v_column_2/res0_in vdd b2b b0a b1b b4b rheo_3v_column_1/out_4 b1a b2b b1b
+ vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b vdd b0b
+ rheo_3v_column_2/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b b2a rheo_3v_column_odd
Xrheo_3v_column_odd_2 b5a b6a rheo_3v_column_2/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b6b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_3/out_5 b1b
+ rheo_3v_column_2/dum1_out rheo_3v_column_3/res0_in vdd b2b b0a b1b b4b rheo_3v_column_2/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_3/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_3 b5a vdd rheo_3v_column_3/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_3/in_5 b0a b3b b0a b0b b3a b1b vss b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_odd_3/in_5
+ b1b rheo_3v_column_3/dum1_out rheo_3v_column_4/res0_in vdd b2b b0a b1b b4b rheo_3v_column_3/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_4/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_4 b5a b6b rheo_3v_column_4/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b6a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_5/out_5 b1b
+ rheo_3v_column_4/dum1_out rheo_3v_column_5/res0_in vdd b2b b0a b1b b4b rheo_3v_column_4/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_5/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_5 b5a b7a rheo_3v_column_5/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b7b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b out b1b rheo_3v_column_5/dum1_out
+ rheo_3v_column_6/res0_in vdd b2b b0a b1b b4b rheo_3v_column_5/out_4 b1a b2b b1b
+ vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b vdd b0b
+ rheo_3v_column_6/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b b2a rheo_3v_column_odd
Xrheo_3v_column_odd_6 b5a b6a rheo_3v_column_6/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b6b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_7/out_5 b1b
+ rheo_3v_column_6/dum1_out rheo_3v_column_7/res0_in vdd b2b b0a b1b b4b rheo_3v_column_6/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_7/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_7 b5a vdd rheo_3v_column_7/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_7/in_5 b0a b3b b0a b0b b3a b1b vss b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_odd_7/in_5
+ b1b rheo_3v_column_7/dum1_out Vlow vdd b2b b0a b1b b4b rheo_3v_column_7/out_4 b1a
+ b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b
+ vdd b0b rheo_3v_column_odd_7/dum_out1 b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_dummy_0 b0a b1b b2a b1a b0b vss vdd b0a b0b vss vdd b0b b0a b0a b0b
+ b0a b0b b0b b0a vdd b0b b0a b2b b1a b0b b0a b0b vss vdd b0a vdd vdd vdd vss vdd
+ b0b vdd b0a b0b b4a b0a b0b b1a vdd b0a vdd b0b vdd b1b b0a vdd b2b vss vss b4b
+ vdd b1b b3a b1a b2b b2a b1a vdd b1a b1b vdd b3b b3a b1b b1a b2a b2b b1a b1b b3b
+ b5b vss vss b5a b1b b1b vdd vdd vdd b0a b0b Vhigh b0a b2a m1_6292_841# b0b rheo_3v_column_0/dum0_in
+ b0a b0b m1_6292_841# vss rheo_3v_column_dummy
Xrheo_3v_column_dummy_1 b0a b1b b2a b1a b0b vss vdd b0a b0b vss vdd b0b b0a b0a b0b
+ b0a b0b b0b b0a vdd b0b b0a b2b b1a b0b b0a b0b vss vdd b0a vdd vdd vdd vss vdd
+ b0b vdd b0a b0b b4a b0a b0b b1a vdd b0a vdd b0b vdd b1b b0a vdd b2b vss vss b4b
+ vdd b1b b3a b1a b2b b2a b1a vdd b1a b1b vdd b3b b3a b1b b1a b2a b2b b1a b1b b3b
+ b5b vss vss b5a b1b b1b vdd vdd vdd b0a b0b m1_25337_837# b0a b2a Vlow b0b m1_25337_837#
+ b0a b0b rheo_3v_column_odd_7/dum_out1 vss rheo_3v_column_dummy
Xrheo_level_shifter_array_0 b0 b3b b3a b4 b0a b4a b7a b1 b0b b5 b4b b7b b1b b5a b1a
+ b6 b2 b5b b6b b2b b2a b3 b7 dvdd vdd b6a dvss rheo_level_shifter_array
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6 a_29_n311# a_n129_n311# a_n29_n214# a_n187_n214#
+ a_129_n214# w_n387_n512#
X0 a_129_n214# a_29_n311# a_n29_n214# w_n387_n512# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X1 a_n29_n214# a_n129_n311# a_n187_n214# w_n387_n512# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U62SY6 a_n108_n464# a_n50_n561# w_n308_n762#
+ a_50_n464#
X0 a_50_n464# a_n50_n561# a_n108_n464# w_n308_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQFX__0 a_129_n200# a_29_n288# a_n129_n288#
+ a_n321_n422# a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6NWY6 w_n387_n762# a_29_n561# a_n129_n561# a_n29_n464#
+ a_n187_n464# a_129_n464#
X0 a_129_n464# a_29_n561# a_n29_n464# w_n387_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X1 a_n29_n464# a_n129_n561# a_n187_n464# w_n387_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8__0 a_50_n200# a_n242_n422# a_n108_n200#
+ a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt balanced_switch hold out in vdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6_0 holdb holdb vdd holdp holdp vdd sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6
Xsky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 out holdb vdd out sky130_fd_pr__pfet_g5v0d10v5_U62SY6
Xsky130_fd_pr__pfet_g5v0d10v5_U62SY6_1 in holdb vdd in sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM1 out holdb holdb vss in out sky130_fd_pr__nfet_g5v0d10v5_EJGQFX__0
Xsky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0 vdd holdp holdp in out out sky130_fd_pr__pfet_g5v0d10v5_U6NWY6
XXM3 in vss in holdp sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8__0
XXM5 out vss out holdp sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8__0
XXM7 hold hold vdd holdb holdb vdd sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6
XXM8 holdb vss vss hold sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8__0
XXD1 vss hold sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
XXM10 holdp vss vss holdb sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8__0
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW__0 a_1293_n197# a_n761_n197# a_1235_n100#
+ a_n1551_n197# a_761_n100# a_n29_n100# a_1393_n100# a_1451_n197# a_n187_n100# a_1551_n100#
+ a_n819_n100# a_n345_n100# a_n1609_n100# a_29_n197# a_n977_n100# a_n1135_n100# a_n129_n197#
+ a_187_n197# a_129_n100# a_n503_n100# a_n1293_n100# a_n287_n197# a_819_n197# a_n661_n100#
+ a_345_n197# a_n1077_n197# a_287_n100# a_n1451_n100# a_n919_n197# a_977_n197# a_n445_n197#
+ a_919_n100# a_503_n197# a_n1235_n197# a_445_n100# w_n1809_n397# a_1077_n100# a_1135_n197#
+ a_n603_n197# a_n1393_n197# a_661_n197# a_603_n100#
X0 a_287_n100# a_187_n197# a_129_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_1235_n100# a_1135_n197# a_1077_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_919_n100# a_819_n197# a_761_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_445_n100# a_345_n197# a_287_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_603_n100# a_503_n197# a_445_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n1293_n100# a_n1393_n197# a_n1451_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n1451_n100# a_n1551_n197# a_n1609_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X7 a_n977_n100# a_n1077_n197# a_n1135_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_n1135_n100# a_n1235_n197# a_n1293_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n661_n100# a_n761_n197# a_n819_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_129_n100# a_29_n197# a_n29_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_n187_n100# a_n287_n197# a_n345_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_n819_n100# a_n919_n197# a_n977_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_n345_n100# a_n445_n197# a_n503_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_n503_n100# a_n603_n197# a_n661_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_n29_n100# a_n129_n197# a_n187_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 a_1393_n100# a_1293_n197# a_1235_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 a_1077_n100# a_977_n197# a_919_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_1551_n100# a_1451_n197# a_1393_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X19 a_761_n100# a_661_n197# a_603_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0 a_50_n100# a_n242_n322# a_n108_n100#
+ a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLJMY6__0 a_n208_n197# a_208_n100# a_n50_n197#
+ a_50_n100# a_n108_n100# w_n466_n397# a_n266_n100# a_108_n197#
X0 a_208_n100# a_108_n197# a_50_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_50_n100# a_n50_n197# a_n108_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n108_n100# a_n208_n197# a_n266_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLWMS5__0 a_n29_n100# a_n187_n100# w_n545_n397#
+ a_n345_n100# a_29_n197# a_n129_n197# a_187_n197# a_129_n100# a_n287_n197# a_287_n100#
X0 a_287_n100# a_187_n197# a_129_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_129_n100# a_29_n197# a_n29_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n187_n100# a_n287_n197# a_n345_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n29_n100# a_n129_n197# a_n187_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_HLA228__0 a_131_1150# a_131_n1582# a_n201_n1582#
+ a_n35_n1582# a_n201_1150# a_n35_1150# a_n331_n1712#
X0 a_n35_1150# a_n35_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X1 a_n201_1150# a_n201_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X2 a_131_1150# a_131_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQFC__0 a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y__0 a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_BH6ZTK__0 a_n29_n100# a_209_n100# a_n209_n188#
+ a_n401_n322# a_n267_n100# a_29_n188#
X0 a_n29_n100# a_n209_n188# a_n267_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.9
X1 a_209_n100# a_29_n188# a_n29_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.9
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ__0 a_n345_118# a_1393_n2934# a_977_n851#
+ a_603_n1626# a_n1451_2734# a_1551_n2498# a_29_n415# a_n661_554# a_n1551_21# a_1451_1329#
+ a_445_118# a_n445_n851# a_n129_n2595# a_761_554# a_n129_1765# a_n661_2298# a_n187_n754#
+ a_29_n1287# a_n977_n2062# a_345_893# a_287_2298# a_1235_n1626# a_n129_n415# a_977_n3031#
+ a_n1235_n2595# a_445_1862# a_761_n2498# a_n29_n2498# a_603_n318# a_187_1765# a_n503_1426#
+ a_29_2637# a_n1235_n851# a_129_1426# a_919_2734# a_1077_990# a_n287_457# a_187_n415#
+ a_n603_n2595# a_445_n1626# a_n977_990# a_n1293_1426# a_n603_2201# a_1393_n2498#
+ a_n1451_2298# a_1135_2201# a_977_21# a_503_n851# a_919_n1626# a_n1393_2201# a_n1135_n2934#
+ a_n129_2637# a_29_n2159# a_1077_n1626# a_n1609_n2934# a_661_2201# a_187_21# a_n1077_n2595#
+ a_445_2734# a_n187_118# a_1551_n754# a_n503_n2934# a_29_457# a_187_2637# a_129_990#
+ a_287_118# a_1077_1862# a_503_n2595# a_n819_n754# a_n287_1765# a_n445_n2595# a_287_n1626#
+ a_919_2298# a_1235_n318# a_187_893# a_1451_457# a_n287_n415# a_n919_n2595# a_1551_n1626#
+ a_1135_n2595# a_n1551_n2595# a_1451_21# a_n129_n1723# a_n1135_n2498# a_819_1765#
+ a_n603_n851# a_761_n318# a_1135_n851# a_n661_1426# a_n345_n754# a_n1609_n2498# a_819_n415#
+ a_n1393_n851# a_287_1426# a_445_2298# a_n761_2201# a_n919_457# a_n345_n2934# a_n1077_1765#
+ a_n1609_n754# a_n1235_n1723# a_n503_n2498# a_n1609_990# a_1293_2201# a_761_n1626#
+ a_603_1862# a_1077_2734# a_661_n851# a_n29_n1626# a_345_n2595# a_n1235_893# a_n445_21#
+ a_n819_n2934# a_n1077_n415# a_503_457# a_n287_n2595# a_n287_2637# a_345_1765# a_n1451_n2934#
+ a_819_n2595# a_n603_n1723# a_345_n415# a_1393_n1626# a_n1451_1426# a_n1393_n2595#
+ a_n1135_n754# a_819_2637# a_n819_118# a_n129_n1287# a_n29_n318# a_n1551_2201# a_n29_990#
+ a_1235_554# a_n919_1765# a_n1135_554# a_919_118# a_n977_n754# a_1551_990# a_n761_457#
+ a_n187_n2934# a_1393_n318# a_n1077_n1723# a_n1451_990# a_n1077_2637# a_n345_n2498#
+ a_n761_n2595# a_n919_n415# a_1293_457# a_n1235_n1287# a_819_893# a_603_2734# a_187_n2595#
+ a_1077_2298# a_n819_n2498# a_345_2637# a_977_1765# a_n761_n851# a_503_n1723# a_n1293_n2934#
+ a_1235_1862# a_1451_n2595# a_1293_n851# a_n445_n1723# a_n1451_n2498# a_29_1329#
+ a_n1077_21# a_129_n1190# a_n445_1765# a_n603_n1287# a_919_1426# a_977_n415# a_n503_990#
+ a_n919_n1723# a_n661_118# a_n445_n415# a_n129_n2159# a_n661_n2934# a_1135_n1723#
+ a_761_1862# a_603_990# a_n1551_n1723# a_n1135_n1626# a_n129_1329# a_761_118# a_n919_2637#
+ a_n187_n318# a_n1077_893# a_345_457# a_661_n2595# a_n1609_n1626# a_n187_n2498# a_345_21#
+ a_n1077_n1287# a_661_893# a_29_21# a_n503_n754# a_n1235_n2159# a_n1551_n851# a_445_1426#
+ a_603_2298# a_129_n754# a_n503_n1626# a_n1235_1765# a_603_n1190# a_n1293_n754# a_187_1329#
+ a_1451_2201# a_977_2637# a_345_n1723# a_1293_n2595# a_1235_2734# a_n287_n1723# a_n1293_n2498#
+ a_503_n1287# a_n1235_n415# a_129_n2062# a_n445_n1287# a_n129_893# a_n445_2637# a_n977_554#
+ a_1077_554# a_n603_n2159# a_503_1765# a_819_n1723# a_1393_990# a_1235_n1190# a_n1293_990#
+ a_n919_n1287# a_503_n415# a_n29_1862# a_761_2734# a_n1393_n1723# a_1135_n1287# a_n661_n2498#
+ a_n1551_n1287# a_n977_n2934# a_1393_1862# a_n1077_n2159# a_977_n2595# a_n761_n1723#
+ a_1551_n318# a_n345_n1626# a_445_n1190# a_603_n2062# a_n1235_2637# a_n345_990# a_129_554#
+ a_187_n1723# a_1077_1426# a_345_n1287# a_n603_21# a_n819_n1626# a_503_n2159# a_919_n1190#
+ a_1235_2298# a_445_990# a_n819_n318# a_n287_n1287# a_n287_1329# a_n445_n2159# a_29_n3031#
+ a_503_2637# a_1451_n1723# a_n1451_n1626# a_187_457# a_819_n1287# a_1451_n851# a_1077_n1190#
+ a_1235_n2062# a_n919_n2159# a_n603_1765# a_n661_n754# a_1135_1765# a_n29_2734# a_n1393_n1287#
+ a_1135_n2159# a_761_2298# a_287_n754# a_n1551_n2159# a_819_1329# a_n187_1862# a_n1393_1765#
+ a_n603_n415# a_1135_n415# a_1393_2734# a_n977_n2498# a_n1393_n415# a_n345_n318#
+ a_661_n1723# a_661_1765# a_n187_n1626# a_n1609_n318# a_287_n1190# a_445_n2062# a_n1077_1329#
+ a_n761_n1287# a_n1609_554# a_603_1426# a_187_n1287# a_n1235_457# a_661_n415# a_345_n2159#
+ a_1551_n1190# a_919_n2062# a_n287_n2159# a_n1451_n754# a_345_1329# a_1293_n1723#
+ a_n1551_893# a_n1293_n1626# a_1451_n1287# a_819_n2159# a_1077_n2062# a_n603_2637#
+ a_n1235_21# a_1135_2637# a_n29_2298# a_n1135_n318# a_n1393_n2159# a_n187_2734# a_n1393_2637#
+ a_n187_990# a_n661_n1626# a_761_n1190# a_n29_554# a_1235_118# a_n919_1329# a_1393_2298#
+ a_n1135_118# a_n977_n318# a_n29_n1190# a_287_990# a_661_n1287# a_n603_893# a_661_2637#
+ a_1551_554# a_287_n2062# a_n1451_554# a_1551_1862# a_n761_n2159# a_1135_893# a_503_21#
+ a_977_n1723# a_819_457# a_n761_1765# a_187_n2159# a_1293_1765# a_1393_n1190# a_1551_n2062#
+ a_919_n754# a_n819_1862# a_n761_n415# a_977_1329# a_1293_n1287# a_1235_1426# a_1451_n2159#
+ a_1293_n415# a_n445_1329# a_n503_554# a_n187_2298# a_761_1426# a_603_554# a_761_n2062#
+ a_n1077_457# a_445_n754# a_n29_n2062# a_n345_1862# a_n1551_1765# a_n977_n1626# a_661_n2159#
+ a_n1393_893# a_1551_2734# a_n1609_1862# a_29_2201# a_661_457# a_n1551_n415# a_n503_n318#
+ a_n761_2637# a_977_n1287# a_129_n318# a_1393_n2062# a_1293_2637# a_n1235_1329# a_n819_2734#
+ a_n1293_n318# a_n129_n3031# a_1293_n2159# a_n129_457# a_n129_2201# a_1077_118# a_n819_990#
+ a_n977_118# a_n1135_n1190# a_503_1329# a_n445_893# a_1393_554# a_919_990# a_n1135_1862#
+ a_n1293_554# a_1135_21# a_n1609_n1190# a_n1235_n3031# a_n29_1426# a_n919_21# a_n345_2734#
+ a_n1551_2637# a_n503_n1190# a_977_893# a_n977_1862# a_187_2201# a_1393_1426# a_n1609_2734#
+ a_1551_2298# a_1077_n754# a_n761_21# a_977_n2159# a_n603_n3031# a_n129_21# a_n345_554#
+ a_129_118# a_n819_2298# a_29_n851# a_1451_1765# a_n661_990# a_445_554# a_n1135_n2062#
+ a_129_n2934# a_761_990# a_1451_n415# a_n1135_2734# a_n1077_n3031# a_n603_1329# a_n661_n318#
+ a_n1609_n2062# a_1135_1329# a_n129_n851# a_287_n318# a_n187_1426# a_n1393_1329#
+ a_n345_n1190# a_n503_n2062# a_n977_2734# a_n345_2298# a_503_n3031# a_603_n754# a_n1609_2298#
+ a_n287_2201# a_n819_n1190# a_n445_n3031# a_n503_1862# a_661_1329# a_129_1862# a_n1609_118#
+ a_n1451_n1190# a_187_n851# a_n287_893# a_603_n2934# a_n1293_1862# a_n919_n3031#
+ a_n1393_21# a_1451_2637# a_1135_n3031# a_n1551_n3031# a_n1451_n318# a_819_2201#
+ a_n1551_457# a_129_n2498# a_29_n2595# a_n1135_2298# a_1235_n2934# a_819_21# a_n1077_2201#
+ a_n187_n1190# a_n345_n2062# a_n187_554# a_n977_2298# a_661_21# w_n1809_n3231# a_n29_118#
+ a_345_n3031# a_29_893# a_n819_n2062# a_n287_n3031# a_n503_2734# a_n603_457# a_287_554#
+ a_345_2201# a_1551_118# a_n1451_118# a_1551_1426# a_129_2734# a_n1293_n1190# a_819_n3031#
+ a_1135_457# a_n1451_n2062# a_445_n2934# a_n1293_2734# a_1235_n754# a_n761_1329#
+ a_603_n2498# a_1451_893# a_1293_1329# a_919_n318# a_n287_n851# a_n1393_n3031# a_n819_1426#
+ a_919_n2934# a_n661_n1190# a_n919_2201# a_761_n754# a_1077_n2934# a_n661_1862# a_1235_n2498#
+ a_n503_118# a_819_n851# a_287_1862# a_n761_n3031# a_n187_n2062# a_603_118# a_187_n3031#
+ a_n919_893# a_445_n318# a_n345_1426# a_n1551_1329# a_n503_2298# a_977_2201# a_n1393_457#
+ a_n1077_n851# a_1451_n3031# a_503_893# a_n1609_1426# a_n1293_n2062# a_287_n2934#
+ a_129_2298# a_n445_2201# a_445_n2498# a_n1293_2298# a_345_n851# a_1551_n2934# a_n1451_1862#
+ a_919_n2498# a_1293_21# a_n819_554# a_n661_n2062# a_n29_n754# a_129_n1626# a_n661_2734#
+ a_29_n1723# a_661_n3031# a_1077_n2498# a_1235_990# a_n445_457# a_919_554# a_1393_118#
+ a_n1135_990# a_n977_n1190# a_n1135_1426# a_287_2734# a_n1293_118# a_n761_893# a_1393_n754#
+ a_n919_n851# a_761_n2934# a_1293_893# a_n1235_2201# a_977_457# a_n977_1426# a_n29_n2934#
+ a_n287_21# a_1293_n3031# a_1077_n318# a_287_n2498# a_503_2201# a_29_1765# a_919_1862#
X0 a_n1135_n318# a_n1235_n415# a_n1293_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_1235_2298# a_1135_2201# a_1077_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_761_554# a_661_457# a_603_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n1135_2298# a_n1235_2201# a_n1293_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n29_990# a_n129_893# a_n187_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_603_118# a_503_21# a_445_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_445_n2498# a_345_n2595# a_287_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_1077_n1626# a_977_n1723# a_919_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_919_n2934# a_819_n3031# a_761_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n1451_n1626# a_n1551_n1723# a_n1609_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X10 a_919_n1190# a_819_n1287# a_761_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_1393_990# a_1293_893# a_1235_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_287_554# a_187_457# a_129_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_129_n2062# a_29_n2159# a_n29_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_n29_n754# a_n129_n851# a_n187_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_603_n754# a_503_n851# a_445_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 a_n1135_1862# a_n1235_1765# a_n1293_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 a_1235_1862# a_1135_1765# a_1077_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_1235_554# a_1135_457# a_1077_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X19 a_1077_n2934# a_977_n3031# a_919_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 a_n1451_n1190# a_n1551_n1287# a_n1609_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X21 a_n1451_n2934# a_n1551_n3031# a_n1609_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X22 a_919_n2498# a_819_n2595# a_761_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 a_1077_n1190# a_977_n1287# a_919_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 a_1077_990# a_977_893# a_919_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 a_919_554# a_819_457# a_761_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 a_n345_n1626# a_n445_n1723# a_n503_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X27 a_445_554# a_345_457# a_287_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X28 a_1551_990# a_1451_893# a_1393_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X29 a_n1293_118# a_n1393_21# a_n1451_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 a_445_n2062# a_345_n2159# a_287_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 a_n819_1426# a_n919_1329# a_n977_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 a_1077_n2498# a_977_n2595# a_919_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 a_n1451_n2498# a_n1551_n2595# a_n1609_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X34 a_n345_n2934# a_n445_n3031# a_n503_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 a_n345_n1190# a_n445_n1287# a_n503_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X36 a_1235_n754# a_1135_n851# a_1077_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 a_n661_1426# a_n761_1329# a_n819_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 a_n1135_n754# a_n1235_n851# a_n1293_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X39 a_761_990# a_661_893# a_603_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 a_n819_n1626# a_n919_n1723# a_n977_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 a_n819_2734# a_n919_2637# a_n977_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X42 a_603_554# a_503_457# a_445_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 a_n1451_118# a_n1551_21# a_n1609_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X44 a_n977_n1626# a_n1077_n1723# a_n1135_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X45 a_n345_n2498# a_n445_n2595# a_n503_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 a_919_n2062# a_819_n2159# a_761_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X47 a_919_1426# a_819_1329# a_761_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X48 a_n661_2734# a_n761_2637# a_n819_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 a_n819_n2934# a_n919_n3031# a_n977_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X50 a_1235_n1626# a_1135_n1723# a_1077_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X51 a_287_990# a_187_893# a_129_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X52 a_n819_n318# a_n919_n415# a_n977_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X53 a_n819_n1190# a_n919_n1287# a_n977_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X54 a_n819_2298# a_n919_2201# a_n977_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X55 a_1235_990# a_1135_893# a_1077_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X56 a_n977_118# a_n1077_21# a_n1135_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 a_n187_1426# a_n287_1329# a_n345_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 a_761_1426# a_661_1329# a_603_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X59 a_n977_n2934# a_n1077_n3031# a_n1135_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X60 a_1077_n2062# a_977_n2159# a_919_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X61 a_n1451_n2062# a_n1551_n2159# a_n1609_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X62 a_n977_n1190# a_n1077_n1287# a_n1135_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X63 a_919_2734# a_819_2637# a_761_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X64 a_n661_n318# a_n761_n415# a_n819_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X65 a_1393_n1626# a_1293_n1723# a_1235_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X66 a_919_990# a_819_893# a_761_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X67 a_1235_n2934# a_1135_n3031# a_1077_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X68 a_n661_2298# a_n761_2201# a_n819_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X69 a_n819_n2498# a_n919_n2595# a_n977_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X70 a_603_n1626# a_503_n1723# a_445_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X71 a_1235_n1190# a_1135_n1287# a_1077_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X72 a_445_990# a_345_893# a_287_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X73 a_761_2734# a_661_2637# a_603_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X74 a_n1293_554# a_n1393_457# a_n1451_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X75 a_n187_2734# a_n287_2637# a_n345_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X76 a_n1135_118# a_n1235_21# a_n1293_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X77 a_919_n318# a_819_n415# a_761_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X78 a_n977_n2498# a_n1077_n2595# a_n1135_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X79 a_n819_1862# a_n919_1765# a_n977_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X80 a_919_2298# a_819_2201# a_761_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X81 a_1393_n2934# a_1293_n3031# a_1235_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X82 a_n345_n2062# a_n445_n2159# a_n503_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X83 a_287_1426# a_187_1329# a_129_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X84 a_1235_n2498# a_1135_n2595# a_1077_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X85 a_761_n1626# a_661_n1723# a_603_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X86 a_1393_n1190# a_1293_n1287# a_1235_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X87 a_603_n2934# a_503_n3031# a_445_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X88 a_n661_1862# a_n761_1765# a_n819_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X89 a_n187_n318# a_n287_n415# a_n345_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X90 a_761_n318# a_661_n415# a_603_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X91 a_603_n1190# a_503_n1287# a_445_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X92 a_1393_1426# a_1293_1329# a_1235_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X93 a_n187_2298# a_n287_2201# a_n345_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X94 a_761_2298# a_661_2201# a_603_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X95 a_n1293_1426# a_n1393_1329# a_n1451_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X96 a_603_990# a_503_893# a_445_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X97 a_n1451_554# a_n1551_457# a_n1609_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X98 a_287_2734# a_187_2637# a_129_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X99 a_761_n2934# a_661_n3031# a_603_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X100 a_1393_n2498# a_1293_n2595# a_1235_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X101 a_919_1862# a_819_1765# a_761_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X102 a_603_n2498# a_503_n2595# a_445_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X103 a_761_n1190# a_661_n1287# a_603_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X104 a_n661_118# a_n761_21# a_n819_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X105 a_n819_n2062# a_n919_n2159# a_n977_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X106 a_n1293_2734# a_n1393_2637# a_n1451_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X107 a_1393_2734# a_1293_2637# a_1235_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X108 a_n819_n754# a_n919_n851# a_n977_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X109 a_129_118# a_29_21# a_n29_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X110 a_n977_554# a_n1077_457# a_n1135_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X111 a_n187_1862# a_n287_1765# a_n345_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X112 a_761_1862# a_661_1765# a_603_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X113 a_287_n318# a_187_n415# a_129_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X114 a_n977_n2062# a_n1077_n2159# a_n1135_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X115 a_287_2298# a_187_2201# a_129_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X116 a_n661_n754# a_n761_n851# a_n819_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X117 a_761_n2498# a_661_n2595# a_603_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X118 a_1235_n2062# a_1135_n2159# a_1077_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X119 a_n187_118# a_n287_21# a_n345_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X120 a_n1293_n318# a_n1393_n415# a_n1451_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X121 a_1393_n318# a_1293_n415# a_1235_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X122 a_n1293_2298# a_n1393_2201# a_n1451_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X123 a_1393_2298# a_1293_2201# a_1235_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X124 a_n345_1426# a_n445_1329# a_n503_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X125 a_n1293_990# a_n1393_893# a_n1451_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X126 a_n503_n1626# a_n603_n1723# a_n661_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X127 a_n1135_554# a_n1235_457# a_n1293_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X128 a_919_n754# a_819_n851# a_761_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X129 a_n819_118# a_n919_21# a_n977_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X130 a_1393_n2062# a_1293_n2159# a_1235_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X131 a_287_n1626# a_187_n1723# a_129_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X132 a_287_1862# a_187_1765# a_129_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X133 a_603_n2062# a_503_n2159# a_445_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X134 a_129_1426# a_29_1329# a_n29_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X135 a_n345_118# a_n445_21# a_n503_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X136 a_n345_2734# a_n445_2637# a_n503_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X137 a_n187_n754# a_n287_n851# a_n345_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X138 a_761_n754# a_661_n851# a_603_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X139 a_1393_1862# a_1293_1765# a_1235_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X140 a_n503_n2934# a_n603_n3031# a_n661_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X141 a_n661_n1626# a_n761_n1723# a_n819_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X142 a_n1293_1862# a_n1393_1765# a_n1451_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X143 a_n503_n1190# a_n603_n1287# a_n661_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X144 a_n1451_990# a_n1551_893# a_n1609_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X145 a_445_1426# a_345_1329# a_287_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X146 a_287_n2934# a_187_n3031# a_129_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X147 a_761_n2062# a_661_n2159# a_603_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X148 a_287_n1190# a_187_n1287# a_129_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X149 a_129_2734# a_29_2637# a_n29_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X150 a_n345_n318# a_n445_n415# a_n503_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X151 a_n1451_1426# a_n1551_1329# a_n1609_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X152 a_1551_1426# a_1451_1329# a_1393_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X153 a_n661_554# a_n761_457# a_n819_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X154 a_n661_n2934# a_n761_n3031# a_n819_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X155 a_n345_2298# a_n445_2201# a_n503_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X156 a_n503_118# a_n603_21# a_n661_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X157 a_n1135_n1626# a_n1235_n1723# a_n1293_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X158 a_n661_n1190# a_n761_n1287# a_n819_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X159 a_129_554# a_29_457# a_n29_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X160 a_n503_n2498# a_n603_n2595# a_n661_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X161 a_445_2734# a_345_2637# a_287_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X162 a_n977_990# a_n1077_893# a_n1135_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X163 a_287_n754# a_187_n851# a_129_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X164 a_129_n318# a_29_n415# a_n29_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X165 a_287_n2498# a_187_n2595# a_129_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X166 a_1551_2734# a_1451_2637# a_1393_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X167 a_n1451_2734# a_n1551_2637# a_n1609_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X168 a_129_2298# a_29_2201# a_n29_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X169 a_n187_554# a_n287_457# a_n345_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X170 a_n1293_n754# a_n1393_n851# a_n1451_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X171 a_1393_n754# a_1293_n851# a_1235_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X172 a_n1293_n1626# a_n1393_n1723# a_n1451_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X173 a_n29_118# a_n129_21# a_n187_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X174 a_n1135_n1190# a_n1235_n1287# a_n1293_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X175 a_n1135_n2934# a_n1235_n3031# a_n1293_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X176 a_n661_n2498# a_n761_n2595# a_n819_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X177 a_n345_1862# a_n445_1765# a_n503_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X178 a_445_n318# a_345_n415# a_287_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X179 a_1551_n1626# a_1451_n1723# a_1393_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X180 a_n29_n1626# a_n129_n1723# a_n187_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X181 a_445_2298# a_345_2201# a_287_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X182 a_n977_1426# a_n1077_1329# a_n1135_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X183 a_n1135_990# a_n1235_893# a_n1293_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X184 a_1551_n318# a_1451_n415# a_1393_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X185 a_n1451_n318# a_n1551_n415# a_n1609_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X186 a_1551_2298# a_1451_2201# a_1393_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X187 a_1077_1426# a_977_1329# a_919_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X188 a_n819_554# a_n919_457# a_n977_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X189 a_1393_118# a_1293_21# a_1235_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X190 a_n1293_n2934# a_n1393_n3031# a_n1451_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X191 a_n1451_2298# a_n1551_2201# a_n1609_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X192 a_n503_1426# a_n603_1329# a_n661_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X193 a_n345_554# a_n445_457# a_n503_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X194 a_n1293_n1190# a_n1393_n1287# a_n1451_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X195 a_n1135_n2498# a_n1235_n2595# a_n1293_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X196 a_129_1862# a_29_1765# a_n29_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X197 a_n29_n2934# a_n129_n3031# a_n187_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X198 a_n187_n1626# a_n287_n1723# a_n345_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X199 a_n977_2734# a_n1077_2637# a_n1135_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X200 a_1551_n2934# a_1451_n3031# a_1393_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X201 a_n503_n2062# a_n603_n2159# a_n661_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X202 a_n29_n1190# a_n129_n1287# a_n187_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X203 a_1551_n1190# a_1451_n1287# a_1393_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X204 a_1077_118# a_977_21# a_919_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X205 a_1077_2734# a_977_2637# a_919_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X206 a_445_1862# a_345_1765# a_287_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X207 a_287_n2062# a_187_n2159# a_129_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X208 a_n503_2734# a_n603_2637# a_n661_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X209 a_n345_n754# a_n445_n851# a_n503_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X210 a_n1293_n2498# a_n1393_n2595# a_n1451_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X211 a_n1451_1862# a_n1551_1765# a_n1609_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X212 a_1551_1862# a_1451_1765# a_1393_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X213 a_n661_990# a_n761_893# a_n819_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X214 a_1551_118# a_1451_21# a_1393_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X215 a_n977_n318# a_n1077_n415# a_n1135_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X216 a_n187_n2934# a_n287_n3031# a_n345_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X217 a_n661_n2062# a_n761_n2159# a_n819_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X218 a_n503_554# a_n603_457# a_n661_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X219 a_1551_n2498# a_1451_n2595# a_1393_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X220 a_n29_n2498# a_n129_n2595# a_n187_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X221 a_n187_n1190# a_n287_n1287# a_n345_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X222 a_n977_2298# a_n1077_2201# a_n1135_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X223 a_n29_1426# a_n129_1329# a_n187_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X224 a_603_1426# a_503_1329# a_445_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X225 a_129_990# a_29_893# a_n29_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X226 a_1077_n318# a_977_n415# a_919_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X227 a_n503_n318# a_n603_n415# a_n661_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X228 a_1077_2298# a_977_2201# a_919_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X229 a_129_n754# a_29_n851# a_n29_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X230 a_n503_2298# a_n603_2201# a_n661_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X231 a_761_118# a_661_21# a_603_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X232 a_n187_990# a_n287_893# a_n345_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X233 a_n187_n2498# a_n287_n2595# a_n345_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X234 a_n1135_n2062# a_n1235_n2159# a_n1293_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X235 a_n29_554# a_n129_457# a_n187_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X236 a_129_n1626# a_29_n1723# a_n29_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X237 a_n29_2734# a_n129_2637# a_n187_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X238 a_603_2734# a_503_2637# a_445_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X239 a_445_n754# a_345_n851# a_287_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X240 a_n977_1862# a_n1077_1765# a_n1135_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X241 a_1551_n754# a_1451_n851# a_1393_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X242 a_287_118# a_187_21# a_129_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X243 a_n1451_n754# a_n1551_n851# a_n1609_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X244 a_1077_1862# a_977_1765# a_919_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X245 a_n819_990# a_n919_893# a_n977_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X246 a_1393_554# a_1293_457# a_1235_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X247 a_n1293_n2062# a_n1393_n2159# a_n1451_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X248 a_n503_1862# a_n603_1765# a_n661_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X249 a_1235_118# a_1135_21# a_1077_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X250 a_n29_n318# a_n129_n415# a_n187_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X251 a_603_n318# a_503_n415# a_445_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X252 a_129_n2934# a_29_n3031# a_n29_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X253 a_603_2298# a_503_2201# a_445_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X254 a_n1135_1426# a_n1235_1329# a_n1293_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X255 a_1235_1426# a_1135_1329# a_1077_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X256 a_n345_990# a_n445_893# a_n503_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X257 a_1551_n2062# a_1451_n2159# a_1393_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X258 a_n29_n2062# a_n129_n2159# a_n187_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X259 a_129_n1190# a_29_n1287# a_n29_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X260 a_n29_2298# a_n129_2201# a_n187_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X261 a_445_n1626# a_345_n1723# a_287_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X262 a_1077_554# a_977_457# a_919_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X263 a_919_118# a_819_21# a_761_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X264 a_1235_2734# a_1135_2637# a_1077_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X265 a_445_118# a_345_21# a_287_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X266 a_129_n2498# a_29_n2595# a_n29_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X267 a_n187_n2062# a_n287_n2159# a_n345_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X268 a_n1135_2734# a_n1235_2637# a_n1293_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X269 a_1551_554# a_1451_457# a_1393_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X270 a_n977_n754# a_n1077_n851# a_n1135_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X271 a_n503_990# a_n603_893# a_n661_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X272 a_445_n2934# a_345_n3031# a_287_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X273 a_n29_1862# a_n129_1765# a_n187_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X274 a_603_1862# a_503_1765# a_445_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X275 a_445_n1190# a_345_n1287# a_287_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X276 a_1077_n754# a_977_n851# a_919_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X277 a_n503_n754# a_n603_n851# a_n661_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X278 a_919_n1626# a_819_n1723# a_761_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X279 a_1235_n318# a_1135_n415# a_1077_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQFY__0 a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQ24__0 a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt follower_amp__0 vdd out ena in vsub vss
XXM12 m1_651_3930# m1_651_3930# out m1_651_3930# vdd out vdd m1_651_3930# vdd out
+ vdd out out m1_651_3930# out vdd m1_651_3930# m1_651_3930# vdd vdd out m1_651_3930#
+ m1_651_3930# out m1_651_3930# m1_651_3930# out vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ out m1_651_3930# m1_651_3930# vdd vdd vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ m1_651_3930# out sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW__0
XXM13 m1_2399_1244# vss nbias ena sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0
XXM24 pbias vss vss nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0
XXM25 pbias vdd pbias vcomp vdd vdd pbias pbias sky130_fd_pr__pfet_g5v0d10v5_KLJMY6__0
XXM27 vcomp m2_526_2596# vdd vcomp out in out m1_811_2614# in vcomp sky130_fd_pr__pfet_g5v0d10v5_KLWMS5__0
XXM29 m1_811_2614# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0
XXR1 m1_3337_606# vdd m1_604_772# m1_604_772# m1_2399_1244# m1_3337_606# vss sky130_fd_pr__res_xhigh_po_0p35_HLA228__0
XXM1 vss m2_1742_2323# m1_505_3709# m2_1930_2454# out in sky130_fd_pr__nfet_g5v0d10v5_FJGQFC__0
XXM5 vdd m1_505_3709# vdd vdd m2_1930_2454# m2_1930_2454# m2_1930_2454# m2_1930_2454#
+ m2_1930_2454# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5__0
XXXD1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
XXM6 vdd m1_651_3930# vdd vdd m2_3105_2460# m2_3105_2460# m2_3105_2460# m2_3105_2460#
+ m2_3105_2460# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5__0
XXXD2 vss in sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
XXM7 vss vss m2_2845_2323# m2_2845_2323# nbias nbias sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y__0
XXM8 vss vss m2_1742_2323# nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0
XXM9 m2_2845_2323# m2_3105_2460# in vss m1_651_3930# out sky130_fd_pr__nfet_05v0_nvt_BH6ZTK__0
XXM30 m2_526_2596# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS__0
XXM20 out vdd m1_505_3709# out vdd out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd m1_505_3709# out vdd m1_505_3709# out m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd out m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ vdd out vdd m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# out out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# out out out m1_505_3709# m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd out vdd m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out out m1_505_3709# vdd out
+ out out m1_505_3709# vdd vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# out m1_505_3709# vdd m1_505_3709# out
+ m1_505_3709# m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# out vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd out vdd
+ vdd m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# out m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# out out vdd out m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# out out vdd vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709# vdd out vdd out
+ out m1_505_3709# vdd vdd out out out m1_505_3709# m1_505_3709# m1_505_3709# out
+ out vdd out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd vdd out vdd m1_505_3709# vdd
+ out out m1_505_3709# out m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out vdd m1_505_3709#
+ m1_505_3709# vdd out vdd out m1_505_3709# out m1_505_3709# out m1_505_3709# out
+ m1_505_3709# vdd m1_505_3709# out m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd vdd m1_505_3709# m1_505_3709# out vdd vdd vdd
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# out vdd out out m1_505_3709# out out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd out vdd out m1_505_3709# vdd out m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out vdd out vdd
+ out m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# out m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# vdd out out m1_505_3709# vdd vdd out out vdd m1_505_3709#
+ out m1_505_3709# vdd out m1_505_3709# m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out out vdd m1_505_3709#
+ vdd out m1_505_3709# out vdd out m1_505_3709# vdd out out vdd out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# out vdd vdd out vdd out out m1_505_3709# vdd m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# vdd out
+ m1_505_3709# m1_505_3709# out sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ__0
XXM10 nbias vss nbias vss nbias vss vss nbias nbias nbias sky130_fd_pr__nfet_g5v0d10v5_H7BQFY__0
XXM22 m2_526_2596# vss out vss out vss vss m2_526_2596# m2_526_2596# m2_526_2596#
+ sky130_fd_pr__nfet_g5v0d10v5_H7BQ24__0
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_L93GHW a_n162_n162# a_n60_n60#
X0 a_n162_n162# a_n60_n60# sky130_fd_pr__diode_pw2nd_05v5 perim=2.4e+06 area=3.6e+11
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt c1_n550_n500# m3_n650_n600#
X0 c1_n550_n500# m3_n650_n600# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_VCAE9S c2_n751_n500# m4_n851_n600#
X0 c2_n751_n500# m4_n851_n600# sky130_fd_pr__cap_mim_m3_2 l=5 w=5
.ends

.subckt hold_cap_array holdval vss
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt
XXC2[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
.ends

.subckt sky130_ef_ip__samplehold out vdd hold in dvdd ena vss dvss
Xx1 x1/hold x3/in x1/in vdd vss balanced_switch
Xx3 vdd out x3/ena x3/in dvss vss follower_amp__0
Xx2 vdd x1/in x3/ena in dvss vss follower_amp__0
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 ena dvdd dvss vdd vdd x3/ena vdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_1 hold dvdd dvss vdd vdd x1/hold vdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 dvss hold sky130_fd_pr__diode_pw2nd_05v5_L93GHW
Xsky130_fd_pr__diode_pw2nd_05v5_L93GHW_1 dvss ena sky130_fd_pr__diode_pw2nd_05v5_L93GHW
Xhold_cap_array_0 x3/in vss hold_cap_array
.ends

.subckt sky130_fd_pr__nfet_01v8_PVEW3M a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_XPB8Y6 a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt Stage0_clk_inv dvddb clka clk clkb dvss
XXM6 dvss clkb dvss clk sky130_fd_pr__nfet_01v8_PVEW3M
XXM8 clkb clka dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
XXM21 dvss clka dvss clkb sky130_fd_pr__nfet_01v8_PVEW3M
XXM22 clk clkb dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8_hvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_03v3_nvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_3HY9VM w_n296_n419# a_n100_n297# a_100_n200# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n296_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt Stage2_latch dvdd enab clkb vout oneg opos dvddb dvss
XXM12 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM15 dvss dvss m2_1568_n2406# clkb sky130_fd_pr__nfet_03v3_nvt_WSEQJ8
XXM18 dvss dvss vout m1_683_n2348# sky130_fd_pr__nfet_01v8_PVEW3M
XXM19 dvddb m1_683_n2348# dvddb vout sky130_fd_pr__pfet_01v8_3HY9VM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_0 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM1 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_1 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_3 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_2 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM2 dvss m1_1866_n2368# m1_683_n2348# opos sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_4 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM3 dvss m2_1568_n2406# m1_1866_n2368# m2_1331_n391# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_5 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM4 dvss m1_2747_n2368# m2_1331_n391# oneg sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM5 dvss m2_1568_n2406# m1_2747_n2368# m1_683_n2348# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM10 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM11 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGL9FS a_29_n597# a_n287_n500# a_n229_n597# a_287_n597#
+ a_229_n500# w_n745_n797# a_n545_n500# a_n487_n597# a_n29_n500# a_487_n500#
X0 a_487_n500# a_287_n597# a_229_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_229_n500# a_29_n597# a_n29_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n597# a_n287_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E2TVSU a_1261_n500# a_n1319_n500# a_29_n597#
+ a_n287_n500# a_n1061_n500# a_n745_n597# a_803_n597# a_745_n500# a_n229_n597# a_287_n597#
+ a_n1003_n597# a_229_n500# w_n1519_n797# a_n545_n500# a_1061_n597# a_1003_n500# a_n487_n597#
+ a_n1261_n597# a_n29_n500# a_545_n597# a_487_n500# a_n803_n500#
X0 a_n1061_n500# a_n1261_n597# a_n1319_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X1 a_1003_n500# a_803_n597# a_745_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_487_n500# a_287_n597# a_229_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_745_n500# a_545_n597# a_487_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1261_n500# a_1061_n597# a_1003_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_229_n500# a_29_n597# a_n29_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n29_n500# a_n229_n597# a_n287_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n500# a_n745_n597# a_n803_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_n803_n500# a_n1003_n597# a_n1061_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n287_n500# a_n487_n597# a_n545_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_03v3_nvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt Stage1 avdd clka vinn vinp oneg opos avss dvdd w_608_n4573# dvss enab
Xx1 clka dvdd dvss avdd avdd x1/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xx2 enab dvdd dvss avdd avdd x2/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
XXM3_2 vinp oneg vinp vinp oneg li_n3_908# li_n3_908# vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM1_1 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM1_2 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM5 opos w_608_n4573# w_608_n4573# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM6_1 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM6_2 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM8 oneg w_608_n4573# w_608_n4573# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM4_2 avss avss w_608_n4573# w_608_n4573# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_0 vinp oneg vinp vinp oneg li_n3_908# li_n3_908#
+ vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_1 vinn opos vinn vinn opos li_n3_908# li_n3_908#
+ vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM2_2 vinn opos vinn vinn opos li_n3_908# li_n3_908# vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__nfet_03v3_nvt_FJGQ2Y_0 avss avss w_608_n4573# w_608_n4573# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
.ends

.subckt Stage0_ena_inv dvdd ena enab dvss
XXM24 dvss enab dvss ena sky130_fd_pr__nfet_01v8_PVEW3M
XXM25 ena enab dvdd dvdd sky130_fd_pr__pfet_01v8_XPB8Y6
.ends

.subckt sky130_icrg_ip__ulpcomp2 ena vout vinn vinp clk dvdd avdd avss w_288_n7621#
+ dvss
Xx1 x3/dvddb x2/clka clk x3/clkb dvss Stage0_clk_inv
Xx3 dvdd x4/enab x3/clkb vout x3/oneg x3/opos x3/dvddb dvss Stage2_latch
Xx2 avdd x2/clka vinn vinp x3/oneg x3/opos avss dvdd w_288_n7621# dvss x4/enab Stage1
Xx4 dvdd ena x4/enab dvss Stage0_ena_inv
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLHCT5 a_n345_n200# a_29_n297# a_n129_n297# a_187_n297#
+ a_129_n200# a_n287_n297# a_287_n200# a_n29_n200# a_n187_n200# w_n545_n497#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n297# a_n29_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n297# a_n187_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KL97Y6 a_29_n297# a_n129_n297# a_129_n200# a_n29_n200#
+ w_n387_n497# a_n187_n200#
X0 a_129_n200# a_29_n297# a_n29_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n297# a_n187_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQFX a_129_n200# a_29_n288# a_n129_n288# a_n321_n422#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt simple_analog_switch on off out vdd vss in
XXM12 out off off off in off out out in vdd sky130_fd_pr__pfet_g5v0d10v5_KLHCT5
XXM14 on on out out vdd out sky130_fd_pr__pfet_g5v0d10v5_KL97Y6
XXM16 on on in in vdd in sky130_fd_pr__pfet_g5v0d10v5_KL97Y6
XXM1 out on on vss in out sky130_fd_pr__nfet_g5v0d10v5_EJGQFX
XXM3 out vss out off sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXM5 in vss in off sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
.ends

.subckt simple_analog_switch_ena1v8 dvdd on out avss avdd dvss in
Xsky130_fd_sc_hvl__inv_2_0 simple_analog_switch_0/off dvss dvss avdd avdd simple_analog_switch_0/on
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 sky130_fd_sc_hvl__inv_2_1/A dvss dvss avdd avdd simple_analog_switch_0/off
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 on dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsimple_analog_switch_0 simple_analog_switch_0/on simple_analog_switch_0/off out avdd
+ avss in simple_analog_switch
Xsky130_fd_sc_hvl__decap_4_0 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_1 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SF7DK5 a_n242_n281# a_n108_n50# a_50_n50# a_n50_n147#
X0 a_50_n50# a_n50_n147# a_n108_n50# a_n242_n281# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VDJU7P a_n29_n50# a_n187_n50# a_n321_n281# a_29_n147#
+ a_n129_n147# a_129_n50#
X0 a_129_n50# a_29_n147# a_n29_n50# a_n321_n281# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n147# a_n187_n50# a_n321_n281# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt minimum_analog_switch on off in vdd vss out
XXM1 vss in in off sky130_fd_pr__nfet_g5v0d10v5_SF7DK5
XXM2 vss out out off sky130_fd_pr__nfet_g5v0d10v5_SF7DK5
XXM3 in out vss on on out sky130_fd_pr__nfet_g5v0d10v5_VDJU7P
.ends

.subckt minimal_n_switch_ena1v8 in dvdd on out avdd avss dvss
Xminimum_analog_switch_0 minimum_analog_switch_0/on sky130_fd_sc_hvl__inv_2_1/Y in
+ avdd avss out minimum_analog_switch
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_1/Y dvss dvss avdd avdd minimum_analog_switch_0/on
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 sky130_fd_sc_hvl__inv_2_1/A dvss dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 on dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_0 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt EF_SW_RST VP2 VP1 RST AVSS DVDD DVSS AVDD
Xsimple_analog_switch_ena1v8_1 DVDD RST VP2 AVSS AVDD DVSS AVSS simple_analog_switch_ena1v8
Xminimal_n_switch_ena1v8_0 VP1 DVDD RST AVSS AVDD AVSS DVSS minimal_n_switch_ena1v8
.ends

.subckt EF_AMUX21x sel b vdd1p8 vo a vdd3p3 vss dvss
Xsky130_fd_sc_hd__inv_2_0 sel dvss dvss vdd1p8 vdd1p8 sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2
Xsimple_analog_switch_ena1v8_1 vdd1p8 sel vo vss vdd3p3 dvss a simple_analog_switch_ena1v8
Xsimple_analog_switch_ena1v8_2 vdd1p8 sky130_fd_sc_hd__inv_2_0/Y vo vss vdd3p3 dvss
+ b simple_analog_switch_ena1v8
.ends

.subckt EF_AMUX0201_ARRAY1 SELD2 SELD3 SELD0 D0 SELD1 SELD4 D1 SELD5 SELD9 SELD8 D5
+ SELD7 SELD6 D8 D7 VH VL SELD10 SELD11 D9 D11 D4 DVDD D10 D2 D6 D3 VDD VSS DVSS
Xx1 SELD3 VL DVDD D3 VH VDD VSS DVSS EF_AMUX21x
Xx3 SELD8 VL DVDD D8 VH VDD VSS DVSS EF_AMUX21x
Xx2 SELD4 VL DVDD D4 VH VDD VSS DVSS EF_AMUX21x
Xx4 SELD6 VL DVDD D6 VH VDD VSS DVSS EF_AMUX21x
Xx5 SELD0 VL DVDD D0 VH VDD VSS DVSS EF_AMUX21x
Xx8 SELD2 VL DVDD D2 VH VDD VSS DVSS EF_AMUX21x
Xx9 SELD11 VL DVDD D11 VH VDD VSS DVSS EF_AMUX21x
Xx10 SELD5 VL DVDD D5 VH VDD VSS DVSS EF_AMUX21x
Xx11 SELD1 VL DVDD D1 VH VDD VSS DVSS EF_AMUX21x
Xx12 SELD10 VL DVDD D10 VH VDD VSS DVSS EF_AMUX21x
XEF_AMUX21x_0 SELD9 VL DVDD D9 VH VDD VSS DVSS EF_AMUX21x
XEF_AMUX21x_1 SELD7 VL DVDD D7 VH VDD VSS DVSS EF_AMUX21x
.ends

.subckt cdac_unit_cap m3_80891_n32882# c1_81071_n33152# c2_81071_n33152#
X0 c1_81071_n33152# m3_80891_n32882# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1 c2_81071_n33152# c1_81071_n33152# sky130_fd_pr__cap_mim_m3_2 l=7 w=7
.ends

.subckt cap_array_half cdac_unit_cap_1[4|9]/c2_81071_n33152# cdac_unit_cap_1[3|0]/m3_80891_n32882#
+ cdac_unit_cap_1[7|7]/m3_80891_n32882# cdac_unit_cap_1[6|7]/m3_80891_n32882# cdac_unit_cap_1[6|9]/m3_80891_n32882#
+ cdac_unit_cap_1[6|0]/c2_81071_n33152# cdac_unit_cap_1[2|7]/m3_80891_n32882# cdac_unit_cap_1[8|0]/m3_80891_n32882#
+ cdac_unit_cap_1[5|1]/m3_80891_n32882# cdac_unit_cap_1[3|9]/c2_81071_n33152# cdac_unit_cap_1[2|0]/m3_80891_n32882#
+ cdac_unit_cap_1[7|5]/m3_80891_n32882# cdac_unit_cap_1[5|9]/m3_80891_n32882# cdac_unit_cap_1[5|0]/c2_81071_n33152#
+ cdac_unit_cap_1[8|9]/c2_81071_n33152# cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap_1[7|0]/m3_80891_n32882#
+ cdac_unit_cap_1[2|6]/m3_80891_n32882# cdac_unit_cap_1[2|9]/c2_81071_n33152# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap_1[1|0]/m3_80891_n32882# cdac_unit_cap_1[4|9]/m3_80891_n32882# cdac_unit_cap_1[4|0]/c2_81071_n33152#
+ cdac_unit_cap_1[7|9]/c2_81071_n33152# cdac_unit_cap_1[6|0]/m3_80891_n32882# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap_1[4|4]/c1_81071_n33152# cdac_unit_cap_1[1|9]/c2_81071_n33152# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap_1[5|7]/m3_80891_n32882# cdac_unit_cap_1[1|7]/m3_80891_n32882# cdac_unit_cap_1[3|9]/m3_80891_n32882#
+ cdac_unit_cap_1[3|0]/c2_81071_n33152# cdac_unit_cap_1[5|5]/m3_80891_n32882# cdac_unit_cap_1[6|9]/c2_81071_n33152#
+ cdac_unit_cap_1[6|8]/m3_80891_n32882# cdac_unit_cap_1[8|7]/m3_80891_n32882# cdac_unit_cap_1[5|0]/m3_80891_n32882#
+ cdac_unit_cap_1[8|9]/m3_80891_n32882# cdac_unit_cap_1[8|0]/c2_81071_n33152# cdac_unit_cap_1[2|9]/m3_80891_n32882#
+ cdac_unit_cap_1[2|0]/c2_81071_n33152# cdac_unit_cap_1[5|9]/c2_81071_n33152# caparray_connect_none_8/m3_85388_n19067#
+ cdac_unit_cap_1[4|8]/m3_80891_n32882# cdac_unit_cap_1[4|0]/m3_80891_n32882# cdac_unit_cap_1[7|9]/m3_80891_n32882#
+ cdac_unit_cap_1[7|0]/c2_81071_n33152# cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_99908_n7967#
+ m4_81638_n9537# cdac_unit_cap_1[1|9]/m3_80891_n32882# cdac_unit_cap_1[1|0]/c2_81071_n33152#
+ cdac_unit_cap_1[4|7]/m3_80891_n32882#
Xcdac_unit_cap_1[0|0] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|0] cdac_unit_cap_1[1|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[1|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|0] cdac_unit_cap_1[2|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[2|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|0] cdac_unit_cap_1[3|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[3|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|0] cdac_unit_cap_1[4|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[4|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|0] cdac_unit_cap_1[5|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[5|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|0] cdac_unit_cap_1[6|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[6|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|0] cdac_unit_cap_1[7|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[7|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|0] cdac_unit_cap_1[8|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[8|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|1] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|1] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|1] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|1] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|1] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|1] cdac_unit_cap_1[5|1]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|1]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|1] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|1] cdac_unit_cap_1[7|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|1] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|2] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|2] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|2] cdac_unit_cap_1[2|6]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|6]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|2] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|2] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|2] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|2] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|2] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|2] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|3] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|3] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|3] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|3] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|3] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|3] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|3] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|3] cdac_unit_cap_1[7|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|3] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|4] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|4] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|4] cdac_unit_cap_1[2|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|4] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|4] cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap_1[4|4]/c1_81071_n33152#
+ cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap
Xcdac_unit_cap_1[5|4] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|4] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|4] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|4] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|5] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|5] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|5] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|5] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|5] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|5] cdac_unit_cap_1[5|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|5] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|5] cdac_unit_cap_1[7|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|5] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|6] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|6] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|6] cdac_unit_cap_1[2|6]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|6]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|6] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|6] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|6] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|6] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|6] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|6] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|7] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|7] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|7] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|7] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|7] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|7] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|7] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|7] cdac_unit_cap_1[7|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|7] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|8] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|8] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|8] cdac_unit_cap_1[2|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|8] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|8] cdac_unit_cap_1[4|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|8] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|8] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|8] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|8] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|9] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|9] cdac_unit_cap_1[1|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[1|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|9] cdac_unit_cap_1[2|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[2|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|9] cdac_unit_cap_1[3|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[3|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|9] cdac_unit_cap_1[4|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[4|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|9] cdac_unit_cap_1[5|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[5|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|9] cdac_unit_cap_1[6|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[6|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|9] cdac_unit_cap_1[7|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[7|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|9] cdac_unit_cap_1[8|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[8|9]/c2_81071_n33152#
+ cdac_unit_cap
.ends

.subckt cdac_ratioed_cap c1_81071_n33170# m3_80891_n32900# c2_81071_n33170#
X0 c1_81071_n33170# m3_80891_n32900# sky130_fd_pr__cap_mim_m3_1 l=7.055 w=7
X1 c2_81071_n33170# c1_81071_n33170# sky130_fd_pr__cap_mim_m3_2 l=7.055 w=7
.ends

.subckt EF_BANK_CAP_12 D8 D0 D4 VP1 D9 D5 D1 D2 D6 VSS D7 D3 D10 D11 w_58549_n26640#
+ VP2
Xcap_array_half_0 VSS VSS D8 D11 VSS VSS D11 VSS D7 VSS VSS D9 VSS VSS VSS VSS VSS
+ D8 VSS D9 VSS VSS VSS VSS VSS D10 VSS VSS D10 D9 D10 VSS VSS D6 VSS D10 D11 VSS
+ VSS VSS VSS VSS VSS VP2 D7 VSS VSS VSS VSS VP2 VSS VSS VSS D11 cap_array_half
Xcap_array_half_1 VSS VSS D2 D5 VSS VSS D5 VSS D1 VSS VSS D3 VSS VSS VSS VSS VSS D2
+ VSS D3 VSS VSS VSS VSS VSS D4 VP1 VSS D4 D3 D4 VSS VSS D0 VSS D4 D5 VSS VSS VSS
+ VSS VSS VSS VP1 D1 VSS VSS VSS VSS VP1 VSS VSS VSS D5 cap_array_half
Xcdac_ratioed_cap_0[0] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[1] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[2] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[3] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[4] VP1 VP2 VP2 cdac_ratioed_cap
Xcdac_ratioed_cap_0[5] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[6] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[7] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[8] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[9] VSS VSS VSS cdac_ratioed_cap
.ends

.subckt sky130_ef_ip__cdac3v_12bit SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8 SELD9
+ VDD DVDD OUT RST SELD10 SELD11 OUTNC SELD0 SELD1 VL VH DVSS VSS
Xx1 OUT OUTNC RST VSS DVDD DVSS VDD EF_SW_RST
Xx3 SELD2 SELD3 SELD0 x4/D0 SELD1 SELD4 x4/D1 SELD5 SELD9 SELD8 x4/D5 SELD7 SELD6
+ x4/D8 x4/D7 VH VL SELD10 SELD11 x4/D9 x4/D11 x4/D4 DVDD x4/D10 x4/D2 x4/D6 x4/D3
+ VDD VSS DVSS EF_AMUX0201_ARRAY1
Xx4 x4/D8 x4/D0 x4/D4 OUTNC x4/D9 x4/D5 x4/D1 x4/D2 x4/D6 VSS x4/D7 x4/D3 x4/D10 x4/D11
+ VDD OUT EF_BANK_CAP_12
.ends

.subckt sky130_fd_pr__res_high_po_0p35_AW5QUD a_n35_300# a_n35_n732# VSUBS
X0 a_n35_300# a_n35_n732# VSUBS sky130_fd_pr__res_high_po_0p35 l=3.16
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9992MR a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NHLDUY a_n108_n34# a_n50_n122# a_50_n34# VSUBS
X0 a_50_n34# a_n50_n122# a_n108_n34# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.1885 pd=1.88 as=0.1885 ps=1.88 w=0.65 l=0.5
.ends

.subckt dac_3v_cell m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799# m1_290_1114#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212# m1_663_847# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ m1_300_n125# m1_821_212# m1_814_483# m1_663_212# m1_814_591# w_316_892# m1_814_n125#
+ m1_290_591# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300# m1_155_n223# m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt dac_3v_cell_top m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ w_318_892# m1_290_1114# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212#
+ m1_663_847# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m1_300_n125# m4_97_801#
+ m1_821_212# m4_97_1059# m1_814_483# m1_663_212# m1_814_591# m1_814_n125# m1_290_591#
+ m1_155_n223# m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 m1_824_799# m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt dac_3v_cell_odd m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ m1_290_1114# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212# m1_663_847#
+ m1_155_n223# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m1_300_n125# m1_821_212#
+ m1_814_483# m1_663_212# m1_814_591# w_316_892# m1_814_n125# m1_290_591# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt dac_3v_column_odd m3_31_13582# res_in0 b3_uq0 b0_uq0 b0_uq5 dac_3v_cell_top_0/m4_97_801#
+ b0_uq4 b0_uq11 b2b_uq0 b4 b4b b0b_uq13 b2 b0_uq10 b1_uq5 dac_3v_cell_0[2]/w_316_892#
+ dac_3v_cell_0[1]/w_316_892# b1_uq4 b0 dac_3v_cell_top_0/m4_97_1059# b1_uq6 b0_uq12
+ b0b_uq6 b0b_uq5 m3_30_13212# b0b_uq4 b1_uq0 b0b_uq3 b3b_uq0 b2b_uq2 b0b_uq2 b0b_uq1
+ b0_uq14 b0b_uq14 dac_3v_cell_0[0]/w_316_892# b0b_uq11 b0b_uq0 b0_uq1 b0_uq6 b0b_uq10
+ out_5 b1_uq1 b1 b3b m2_791_14877# m2_801_196# dum_in0 b0b_uq12 b1b_uq6 res_out1
+ b0_uq13 b2_uq2 b2b_uq1 out4 b1b_uq5 dac_3v_cell_0[4]/w_316_892# b2_uq1 b3 dac_3v_cell_odd_0/w_316_892#
+ b1b_uq4 b0_uq3 b2_uq0 b1b_uq3 b1b_uq2 b1b_uq1 b0_uq2 b1_uq2 b1b_uq0 b0b_uq9 m2_791_1314#
+ dac_3v_cell_0[5]/w_316_892# b0_uq9 in_5 b0b dum_out1 b1_uq3 b0_uq8 dac_3v_cell_0[3]/w_316_892#
+ b1b b0b_uq8 b0b_uq7 b0_uq7 m2_801_13759# b2b VSUBS
Xdac_3v_cell_0[0] b0_uq2 dac_3v_cell_odd_0/w_316_892# out0_2 out0_1_0 dac_3v_cell_0[0]/m1_824_799#
+ b2b_uq0 VSUBS out0_0_0 out1_0_3 dac_3v_cell_odd_0/m1_824_799# b0b_uq1 out1_1_1 b1b
+ out1_0_3 b0b_uq2 dac_3v_cell_0[0]/w_316_892# b1 b2_uq0 dac_3v_cell_0[1]/m1_155_n223#
+ dac_3v_cell_0[0]/m1_155_n223# b0_uq1 dac_3v_cell
Xdac_3v_cell_0[1] b0b_uq4 dac_3v_cell_0[0]/w_316_892# out0_0_1 out0_1_0 dac_3v_cell_0[1]/m1_824_799#
+ b1_uq1 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[0]/m1_824_799# b0_uq3 out1_1_1 b2b
+ out1_2 b0_uq4 dac_3v_cell_0[1]/w_316_892# b2 b1b_uq1 dac_3v_cell_0[2]/m1_155_n223#
+ dac_3v_cell_0[1]/m1_155_n223# b0b_uq3 dac_3v_cell
Xdac_3v_cell_0[2] b0_uq6 dac_3v_cell_0[1]/w_316_892# out_3 out0_2 dac_3v_cell_0[2]/m1_824_799#
+ b3b_uq0 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[1]/m1_824_799# b0b_uq5 out1_1_1 b1_uq2
+ out1_0_2 b0b_uq6 dac_3v_cell_0[2]/w_316_892# b1b_uq2 b3_uq0 dac_3v_cell_0[3]/m1_155_n223#
+ dac_3v_cell_0[2]/m1_155_n223# b0_uq5 dac_3v_cell
Xdac_3v_cell_0[3] b0b_uq8 dac_3v_cell_0[2]/w_316_892# out0_0_2 m3_296_8710# dac_3v_cell_0[3]/m1_824_799#
+ b1b_uq3 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[2]/m1_824_799# b0_uq7 out1_2 b3b out_3
+ b0_uq8 dac_3v_cell_0[3]/w_316_892# b3 b1_uq3 dac_3v_cell_0[4]/m1_155_n223# dac_3v_cell_0[3]/m1_155_n223#
+ b0b_uq7 dac_3v_cell
Xdac_3v_cell_0[4] b0_uq10 dac_3v_cell_0[3]/w_316_892# out0_2 m3_296_8710# dac_3v_cell_0[4]/m1_824_799#
+ b2_uq1 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[3]/m1_824_799# b0b_uq9 out1_1_0 b1b_uq4
+ out1_0_1 b0b_uq10 dac_3v_cell_0[4]/w_316_892# b1_uq4 b2b_uq1 dac_3v_cell_0[5]/m1_155_n223#
+ dac_3v_cell_0[4]/m1_155_n223# b0_uq9 dac_3v_cell
Xdac_3v_cell_0[5] b0b_uq12 dac_3v_cell_0[4]/w_316_892# out0_0_3 m3_296_8710# dac_3v_cell_0[5]/m1_824_799#
+ b1_uq5 VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[4]/m1_824_799# b0_uq11 out1_1_0 b2_uq2
+ out1_2 b0_uq12 dac_3v_cell_0[5]/w_316_892# b2b_uq2 b1b_uq5 dac_3v_cell_top_0/m1_155_n223#
+ dac_3v_cell_0[5]/m1_155_n223# b0b_uq11 dac_3v_cell
Xdac_3v_cell_1 m2_791_1314# m2_801_196# m2_329_1119# m2_329_1119# res_out1 m2_791_1314#
+ VSUBS m2_457_485# m2_329_1119# dum_out1 m2_801_196# m2_457_485# VSUBS m2_457_485#
+ VSUBS m2_791_1314# m2_801_196# VSUBS res_in0 dum_in0 VSUBS dac_3v_cell
Xdac_3v_cell_2 m2_791_14877# m2_801_13759# m2_331_14682# m2_331_14682# dum_out0 m2_791_14877#
+ VSUBS m2_458_14048# m2_331_14682# res_in1 m2_801_13759# m2_458_14048# VSUBS m2_458_14048#
+ VSUBS m2_791_14877# m2_801_13759# VSUBS dum_out0 res_in1 VSUBS dac_3v_cell
Xdac_3v_cell_top_0 b0_uq14 dac_3v_cell_0[5]/w_316_892# in_5 out_5 res_in1 m2_801_13759#
+ m3_31_13582# VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[5]/m1_824_799# b0b_uq13 dac_3v_cell_top_0/m4_97_801#
+ out1_1_0 dac_3v_cell_top_0/m4_97_1059# b1_uq6 out1_0_0 b0b_uq14 b1b_uq6 m3_30_13212#
+ dac_3v_cell_top_0/m1_155_n223# b0_uq13 dac_3v_cell_top
Xdac_3v_cell_odd_0 b0b m2_791_1314# out0_0_0 out0_1_0 dac_3v_cell_odd_0/m1_824_799#
+ b1b_uq0 VSUBS out0_0_0 out1_0_3 res_in0 res_out1 b0_uq0 out_3 b4 out4 b0 dac_3v_cell_odd_0/w_316_892#
+ b4b b1_uq0 dac_3v_cell_0[0]/m1_155_n223# b0b_uq0 dac_3v_cell_odd
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW a_1293_n197# a_n761_n197# a_1235_n100#
+ a_n1551_n197# a_761_n100# a_n29_n100# a_1393_n100# a_1451_n197# a_n187_n100# a_1551_n100#
+ a_n819_n100# a_n345_n100# a_n1609_n100# a_29_n197# a_n977_n100# a_n1135_n100# a_n129_n197#
+ a_187_n197# a_129_n100# a_n503_n100# a_n1293_n100# a_n287_n197# a_819_n197# a_n661_n100#
+ a_345_n197# a_n1077_n197# a_287_n100# a_n1451_n100# a_n919_n197# a_977_n197# a_n445_n197#
+ a_919_n100# a_503_n197# a_n1235_n197# a_445_n100# w_n1809_n397# a_1077_n100# a_1135_n197#
+ a_n603_n197# a_n1393_n197# a_661_n197# a_603_n100#
X0 a_287_n100# a_187_n197# a_129_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_1235_n100# a_1135_n197# a_1077_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_919_n100# a_819_n197# a_761_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_445_n100# a_345_n197# a_287_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_603_n100# a_503_n197# a_445_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n1293_n100# a_n1393_n197# a_n1451_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n1451_n100# a_n1551_n197# a_n1609_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X7 a_n977_n100# a_n1077_n197# a_n1135_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_n1135_n100# a_n1235_n197# a_n1293_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n661_n100# a_n761_n197# a_n819_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_129_n100# a_29_n197# a_n29_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_n187_n100# a_n287_n197# a_n345_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_n819_n100# a_n919_n197# a_n977_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_n345_n100# a_n445_n197# a_n503_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_n503_n100# a_n603_n197# a_n661_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_n29_n100# a_n129_n197# a_n187_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 a_1393_n100# a_1293_n197# a_1235_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 a_1077_n100# a_977_n197# a_919_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_1551_n100# a_1451_n197# a_1393_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X19 a_761_n100# a_661_n197# a_603_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQFS a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLJMY6 a_n208_n197# a_208_n100# a_n50_n197# a_50_n100#
+ a_n108_n100# w_n466_n397# a_n266_n100# a_108_n197#
X0 a_208_n100# a_108_n197# a_50_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_50_n100# a_n50_n197# a_n108_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n108_n100# a_n208_n197# a_n266_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLWMS5 a_n29_n100# a_n187_n100# w_n545_n397#
+ a_n345_n100# a_29_n197# a_n129_n197# a_187_n197# a_129_n100# a_n287_n197# a_287_n100#
X0 a_287_n100# a_187_n197# a_129_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_129_n100# a_29_n197# a_n29_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n187_n100# a_n287_n197# a_n345_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n29_n100# a_n129_n197# a_n187_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_HLA228 a_131_1150# a_131_n1582# a_n201_n1582#
+ a_n35_n1582# a_n201_1150# a_n35_1150# a_n331_n1712#
X0 a_n35_1150# a_n35_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X1 a_n201_1150# a_n201_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X2 a_131_1150# a_131_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQFC a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__1 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_BH6ZTK a_n29_n100# a_209_n100# a_n209_n188# a_n401_n322#
+ a_n267_n100# a_29_n188#
X0 a_n29_n100# a_n209_n188# a_n267_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.9
X1 a_209_n100# a_29_n188# a_n29_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.9
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ a_n345_118# a_1393_n2934# a_977_n851#
+ a_603_n1626# a_n1451_2734# a_1551_n2498# a_29_n415# a_n661_554# a_n1551_21# a_1451_1329#
+ a_445_118# a_n445_n851# a_n129_n2595# a_761_554# a_n129_1765# a_n661_2298# a_n187_n754#
+ a_29_n1287# a_n977_n2062# a_345_893# a_287_2298# a_1235_n1626# a_n129_n415# a_977_n3031#
+ a_n1235_n2595# a_445_1862# a_761_n2498# a_n29_n2498# a_603_n318# a_187_1765# a_n503_1426#
+ a_29_2637# a_n1235_n851# a_129_1426# a_919_2734# a_1077_990# a_n287_457# a_187_n415#
+ a_n603_n2595# a_445_n1626# a_n977_990# a_n1293_1426# a_n603_2201# a_1393_n2498#
+ a_n1451_2298# a_1135_2201# a_977_21# a_503_n851# a_919_n1626# a_n1393_2201# a_n1135_n2934#
+ a_n129_2637# a_29_n2159# a_1077_n1626# a_n1609_n2934# a_661_2201# a_187_21# a_n1077_n2595#
+ a_445_2734# a_n187_118# a_1551_n754# a_n503_n2934# a_29_457# a_187_2637# a_129_990#
+ a_287_118# a_1077_1862# a_503_n2595# a_n819_n754# a_n287_1765# a_n445_n2595# a_287_n1626#
+ a_919_2298# a_1235_n318# a_187_893# a_1451_457# a_n287_n415# a_n919_n2595# a_1551_n1626#
+ a_1135_n2595# a_n1551_n2595# a_1451_21# a_n129_n1723# a_n1135_n2498# a_819_1765#
+ a_n603_n851# a_761_n318# a_1135_n851# a_n661_1426# a_n345_n754# a_n1609_n2498# a_819_n415#
+ a_n1393_n851# a_287_1426# a_445_2298# a_n761_2201# a_n919_457# a_n345_n2934# a_n1077_1765#
+ a_n1609_n754# a_n1235_n1723# a_n503_n2498# a_n1609_990# a_1293_2201# a_761_n1626#
+ a_603_1862# a_1077_2734# a_661_n851# a_n29_n1626# a_345_n2595# a_n1235_893# a_n445_21#
+ a_n819_n2934# a_n1077_n415# a_503_457# a_n287_n2595# a_n287_2637# a_345_1765# a_n1451_n2934#
+ a_819_n2595# a_n603_n1723# a_345_n415# a_1393_n1626# a_n1451_1426# a_n1393_n2595#
+ a_n1135_n754# a_819_2637# a_n819_118# a_n129_n1287# a_n29_n318# a_n1551_2201# a_n29_990#
+ a_1235_554# a_n919_1765# a_n1135_554# a_919_118# a_n977_n754# a_1551_990# a_n761_457#
+ a_n187_n2934# a_1393_n318# a_n1077_n1723# a_n1451_990# a_n1077_2637# a_n345_n2498#
+ a_n761_n2595# a_n919_n415# a_1293_457# a_n1235_n1287# a_819_893# a_603_2734# a_187_n2595#
+ a_1077_2298# a_n819_n2498# a_345_2637# a_977_1765# a_n761_n851# a_503_n1723# a_n1293_n2934#
+ a_1235_1862# a_1451_n2595# a_1293_n851# a_n445_n1723# a_n1451_n2498# a_29_1329#
+ a_n1077_21# a_129_n1190# a_n445_1765# a_n603_n1287# a_919_1426# a_977_n415# a_n503_990#
+ a_n919_n1723# a_n661_118# a_n445_n415# a_n129_n2159# a_n661_n2934# a_1135_n1723#
+ a_761_1862# a_603_990# a_n1551_n1723# a_n1135_n1626# a_n129_1329# a_761_118# a_n919_2637#
+ a_n187_n318# a_n1077_893# a_345_457# a_661_n2595# a_n1609_n1626# a_n187_n2498# a_345_21#
+ a_n1077_n1287# a_661_893# a_29_21# a_n503_n754# a_n1235_n2159# a_n1551_n851# a_445_1426#
+ a_603_2298# a_129_n754# a_n503_n1626# a_n1235_1765# a_603_n1190# a_n1293_n754# a_187_1329#
+ a_1451_2201# a_977_2637# a_345_n1723# a_1293_n2595# a_1235_2734# a_n287_n1723# a_n1293_n2498#
+ a_503_n1287# a_n1235_n415# a_129_n2062# a_n445_n1287# a_n129_893# a_n445_2637# a_n977_554#
+ a_1077_554# a_n603_n2159# a_503_1765# a_819_n1723# a_1393_990# a_1235_n1190# a_n1293_990#
+ a_n919_n1287# a_503_n415# a_n29_1862# a_761_2734# a_n1393_n1723# a_1135_n1287# a_n661_n2498#
+ a_n1551_n1287# a_n977_n2934# a_1393_1862# a_n1077_n2159# a_977_n2595# a_n761_n1723#
+ a_1551_n318# a_n345_n1626# a_445_n1190# a_603_n2062# a_n1235_2637# a_n345_990# a_129_554#
+ a_187_n1723# a_1077_1426# a_345_n1287# a_n603_21# a_n819_n1626# a_503_n2159# a_919_n1190#
+ a_1235_2298# a_445_990# a_n819_n318# a_n287_n1287# a_n287_1329# a_n445_n2159# a_29_n3031#
+ a_503_2637# a_1451_n1723# a_n1451_n1626# a_187_457# a_819_n1287# a_1451_n851# a_1077_n1190#
+ a_1235_n2062# a_n919_n2159# a_n603_1765# a_n661_n754# a_1135_1765# a_n29_2734# a_n1393_n1287#
+ a_1135_n2159# a_761_2298# a_287_n754# a_n1551_n2159# a_819_1329# a_n187_1862# a_n1393_1765#
+ a_n603_n415# a_1135_n415# a_1393_2734# a_n977_n2498# a_n1393_n415# a_n345_n318#
+ a_661_n1723# a_661_1765# a_n187_n1626# a_n1609_n318# a_287_n1190# a_445_n2062# a_n1077_1329#
+ a_n761_n1287# a_n1609_554# a_603_1426# a_187_n1287# a_n1235_457# a_661_n415# a_345_n2159#
+ a_1551_n1190# a_919_n2062# a_n287_n2159# a_n1451_n754# a_345_1329# a_1293_n1723#
+ a_n1551_893# a_n1293_n1626# a_1451_n1287# a_819_n2159# a_1077_n2062# a_n603_2637#
+ a_n1235_21# a_1135_2637# a_n29_2298# a_n1135_n318# a_n1393_n2159# a_n187_2734# a_n1393_2637#
+ a_n187_990# a_n661_n1626# a_761_n1190# a_n29_554# a_1235_118# a_n919_1329# a_1393_2298#
+ a_n1135_118# a_n977_n318# a_n29_n1190# a_287_990# a_661_n1287# a_n603_893# a_661_2637#
+ a_1551_554# a_287_n2062# a_n1451_554# a_1551_1862# a_n761_n2159# a_1135_893# a_503_21#
+ a_977_n1723# a_819_457# a_n761_1765# a_187_n2159# a_1293_1765# a_1393_n1190# a_1551_n2062#
+ a_919_n754# a_n819_1862# a_n761_n415# a_977_1329# a_1293_n1287# a_1235_1426# a_1451_n2159#
+ a_1293_n415# a_n445_1329# a_n503_554# a_n187_2298# a_761_1426# a_603_554# a_761_n2062#
+ a_n1077_457# a_445_n754# a_n29_n2062# a_n345_1862# a_n1551_1765# a_n977_n1626# a_661_n2159#
+ a_n1393_893# a_1551_2734# a_n1609_1862# a_29_2201# a_661_457# a_n1551_n415# a_n503_n318#
+ a_n761_2637# a_977_n1287# a_129_n318# a_1393_n2062# a_1293_2637# a_n1235_1329# a_n819_2734#
+ a_n1293_n318# a_n129_n3031# a_1293_n2159# a_n129_457# a_n129_2201# a_1077_118# a_n819_990#
+ a_n977_118# a_n1135_n1190# a_503_1329# a_n445_893# a_1393_554# a_919_990# a_n1135_1862#
+ a_n1293_554# a_1135_21# a_n1609_n1190# a_n1235_n3031# a_n29_1426# a_n919_21# a_n345_2734#
+ a_n1551_2637# a_n503_n1190# a_977_893# a_n977_1862# a_187_2201# a_1393_1426# a_n1609_2734#
+ a_1551_2298# a_1077_n754# a_n761_21# a_977_n2159# a_n603_n3031# a_n129_21# a_n345_554#
+ a_129_118# a_n819_2298# a_29_n851# a_1451_1765# a_n661_990# a_445_554# a_n1135_n2062#
+ a_129_n2934# a_761_990# a_1451_n415# a_n1135_2734# a_n1077_n3031# a_n603_1329# a_n661_n318#
+ a_n1609_n2062# a_1135_1329# a_n129_n851# a_287_n318# a_n187_1426# a_n1393_1329#
+ a_n345_n1190# a_n503_n2062# a_n977_2734# a_n345_2298# a_503_n3031# a_603_n754# a_n1609_2298#
+ a_n287_2201# a_n819_n1190# a_n445_n3031# a_n503_1862# a_661_1329# a_129_1862# a_n1609_118#
+ a_n1451_n1190# a_187_n851# a_n287_893# a_603_n2934# a_n1293_1862# a_n919_n3031#
+ a_n1393_21# a_1451_2637# a_1135_n3031# a_n1551_n3031# a_n1451_n318# a_819_2201#
+ a_n1551_457# a_129_n2498# a_29_n2595# a_n1135_2298# a_1235_n2934# a_819_21# a_n1077_2201#
+ a_n187_n1190# a_n345_n2062# a_n187_554# a_n977_2298# a_661_21# w_n1809_n3231# a_n29_118#
+ a_345_n3031# a_29_893# a_n819_n2062# a_n287_n3031# a_n503_2734# a_n603_457# a_287_554#
+ a_345_2201# a_1551_118# a_n1451_118# a_1551_1426# a_129_2734# a_n1293_n1190# a_819_n3031#
+ a_1135_457# a_n1451_n2062# a_445_n2934# a_n1293_2734# a_1235_n754# a_n761_1329#
+ a_603_n2498# a_1451_893# a_1293_1329# a_919_n318# a_n287_n851# a_n1393_n3031# a_n819_1426#
+ a_919_n2934# a_n661_n1190# a_n919_2201# a_761_n754# a_1077_n2934# a_n661_1862# a_1235_n2498#
+ a_n503_118# a_819_n851# a_287_1862# a_n761_n3031# a_n187_n2062# a_603_118# a_187_n3031#
+ a_n919_893# a_445_n318# a_n345_1426# a_n1551_1329# a_n503_2298# a_977_2201# a_n1393_457#
+ a_n1077_n851# a_1451_n3031# a_503_893# a_n1609_1426# a_n1293_n2062# a_287_n2934#
+ a_129_2298# a_n445_2201# a_445_n2498# a_n1293_2298# a_345_n851# a_1551_n2934# a_n1451_1862#
+ a_919_n2498# a_1293_21# a_n819_554# a_n661_n2062# a_n29_n754# a_129_n1626# a_n661_2734#
+ a_29_n1723# a_661_n3031# a_1077_n2498# a_1235_990# a_n445_457# a_919_554# a_1393_118#
+ a_n1135_990# a_n977_n1190# a_n1135_1426# a_287_2734# a_n1293_118# a_n761_893# a_1393_n754#
+ a_n919_n851# a_761_n2934# a_1293_893# a_n1235_2201# a_977_457# a_n977_1426# a_n29_n2934#
+ a_n287_21# a_1293_n3031# a_1077_n318# a_287_n2498# a_503_2201# a_29_1765# a_919_1862#
X0 a_n1135_n318# a_n1235_n415# a_n1293_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_1235_2298# a_1135_2201# a_1077_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_761_554# a_661_457# a_603_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n1135_2298# a_n1235_2201# a_n1293_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n29_990# a_n129_893# a_n187_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_603_118# a_503_21# a_445_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_445_n2498# a_345_n2595# a_287_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_1077_n1626# a_977_n1723# a_919_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_919_n2934# a_819_n3031# a_761_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n1451_n1626# a_n1551_n1723# a_n1609_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X10 a_919_n1190# a_819_n1287# a_761_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_1393_990# a_1293_893# a_1235_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_287_554# a_187_457# a_129_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_129_n2062# a_29_n2159# a_n29_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_n29_n754# a_n129_n851# a_n187_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_603_n754# a_503_n851# a_445_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 a_n1135_1862# a_n1235_1765# a_n1293_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 a_1235_1862# a_1135_1765# a_1077_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_1235_554# a_1135_457# a_1077_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X19 a_1077_n2934# a_977_n3031# a_919_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 a_n1451_n1190# a_n1551_n1287# a_n1609_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X21 a_n1451_n2934# a_n1551_n3031# a_n1609_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X22 a_919_n2498# a_819_n2595# a_761_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 a_1077_n1190# a_977_n1287# a_919_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 a_1077_990# a_977_893# a_919_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 a_919_554# a_819_457# a_761_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 a_n345_n1626# a_n445_n1723# a_n503_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X27 a_445_554# a_345_457# a_287_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X28 a_1551_990# a_1451_893# a_1393_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X29 a_n1293_118# a_n1393_21# a_n1451_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 a_445_n2062# a_345_n2159# a_287_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 a_n819_1426# a_n919_1329# a_n977_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 a_1077_n2498# a_977_n2595# a_919_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 a_n1451_n2498# a_n1551_n2595# a_n1609_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X34 a_n345_n2934# a_n445_n3031# a_n503_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 a_n345_n1190# a_n445_n1287# a_n503_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X36 a_1235_n754# a_1135_n851# a_1077_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 a_n661_1426# a_n761_1329# a_n819_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 a_n1135_n754# a_n1235_n851# a_n1293_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X39 a_761_990# a_661_893# a_603_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 a_n819_n1626# a_n919_n1723# a_n977_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 a_n819_2734# a_n919_2637# a_n977_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X42 a_603_554# a_503_457# a_445_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 a_n1451_118# a_n1551_21# a_n1609_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X44 a_n977_n1626# a_n1077_n1723# a_n1135_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X45 a_n345_n2498# a_n445_n2595# a_n503_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 a_919_n2062# a_819_n2159# a_761_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X47 a_919_1426# a_819_1329# a_761_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X48 a_n661_2734# a_n761_2637# a_n819_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 a_n819_n2934# a_n919_n3031# a_n977_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X50 a_1235_n1626# a_1135_n1723# a_1077_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X51 a_287_990# a_187_893# a_129_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X52 a_n819_n318# a_n919_n415# a_n977_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X53 a_n819_n1190# a_n919_n1287# a_n977_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X54 a_n819_2298# a_n919_2201# a_n977_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X55 a_1235_990# a_1135_893# a_1077_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X56 a_n977_118# a_n1077_21# a_n1135_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 a_n187_1426# a_n287_1329# a_n345_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 a_761_1426# a_661_1329# a_603_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X59 a_n977_n2934# a_n1077_n3031# a_n1135_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X60 a_1077_n2062# a_977_n2159# a_919_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X61 a_n1451_n2062# a_n1551_n2159# a_n1609_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X62 a_n977_n1190# a_n1077_n1287# a_n1135_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X63 a_919_2734# a_819_2637# a_761_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X64 a_n661_n318# a_n761_n415# a_n819_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X65 a_1393_n1626# a_1293_n1723# a_1235_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X66 a_919_990# a_819_893# a_761_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X67 a_1235_n2934# a_1135_n3031# a_1077_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X68 a_n661_2298# a_n761_2201# a_n819_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X69 a_n819_n2498# a_n919_n2595# a_n977_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X70 a_603_n1626# a_503_n1723# a_445_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X71 a_1235_n1190# a_1135_n1287# a_1077_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X72 a_445_990# a_345_893# a_287_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X73 a_761_2734# a_661_2637# a_603_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X74 a_n1293_554# a_n1393_457# a_n1451_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X75 a_n187_2734# a_n287_2637# a_n345_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X76 a_n1135_118# a_n1235_21# a_n1293_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X77 a_919_n318# a_819_n415# a_761_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X78 a_n977_n2498# a_n1077_n2595# a_n1135_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X79 a_n819_1862# a_n919_1765# a_n977_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X80 a_919_2298# a_819_2201# a_761_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X81 a_1393_n2934# a_1293_n3031# a_1235_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X82 a_n345_n2062# a_n445_n2159# a_n503_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X83 a_287_1426# a_187_1329# a_129_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X84 a_1235_n2498# a_1135_n2595# a_1077_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X85 a_761_n1626# a_661_n1723# a_603_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X86 a_1393_n1190# a_1293_n1287# a_1235_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X87 a_603_n2934# a_503_n3031# a_445_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X88 a_n661_1862# a_n761_1765# a_n819_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X89 a_n187_n318# a_n287_n415# a_n345_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X90 a_761_n318# a_661_n415# a_603_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X91 a_603_n1190# a_503_n1287# a_445_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X92 a_1393_1426# a_1293_1329# a_1235_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X93 a_n187_2298# a_n287_2201# a_n345_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X94 a_761_2298# a_661_2201# a_603_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X95 a_n1293_1426# a_n1393_1329# a_n1451_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X96 a_603_990# a_503_893# a_445_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X97 a_n1451_554# a_n1551_457# a_n1609_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X98 a_287_2734# a_187_2637# a_129_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X99 a_761_n2934# a_661_n3031# a_603_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X100 a_1393_n2498# a_1293_n2595# a_1235_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X101 a_919_1862# a_819_1765# a_761_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X102 a_603_n2498# a_503_n2595# a_445_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X103 a_761_n1190# a_661_n1287# a_603_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X104 a_n661_118# a_n761_21# a_n819_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X105 a_n819_n2062# a_n919_n2159# a_n977_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X106 a_n1293_2734# a_n1393_2637# a_n1451_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X107 a_1393_2734# a_1293_2637# a_1235_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X108 a_n819_n754# a_n919_n851# a_n977_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X109 a_129_118# a_29_21# a_n29_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X110 a_n977_554# a_n1077_457# a_n1135_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X111 a_n187_1862# a_n287_1765# a_n345_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X112 a_761_1862# a_661_1765# a_603_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X113 a_287_n318# a_187_n415# a_129_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X114 a_n977_n2062# a_n1077_n2159# a_n1135_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X115 a_287_2298# a_187_2201# a_129_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X116 a_n661_n754# a_n761_n851# a_n819_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X117 a_761_n2498# a_661_n2595# a_603_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X118 a_1235_n2062# a_1135_n2159# a_1077_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X119 a_n187_118# a_n287_21# a_n345_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X120 a_n1293_n318# a_n1393_n415# a_n1451_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X121 a_1393_n318# a_1293_n415# a_1235_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X122 a_n1293_2298# a_n1393_2201# a_n1451_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X123 a_1393_2298# a_1293_2201# a_1235_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X124 a_n345_1426# a_n445_1329# a_n503_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X125 a_n1293_990# a_n1393_893# a_n1451_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X126 a_n503_n1626# a_n603_n1723# a_n661_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X127 a_n1135_554# a_n1235_457# a_n1293_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X128 a_919_n754# a_819_n851# a_761_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X129 a_n819_118# a_n919_21# a_n977_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X130 a_1393_n2062# a_1293_n2159# a_1235_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X131 a_287_n1626# a_187_n1723# a_129_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X132 a_287_1862# a_187_1765# a_129_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X133 a_603_n2062# a_503_n2159# a_445_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X134 a_129_1426# a_29_1329# a_n29_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X135 a_n345_118# a_n445_21# a_n503_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X136 a_n345_2734# a_n445_2637# a_n503_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X137 a_n187_n754# a_n287_n851# a_n345_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X138 a_761_n754# a_661_n851# a_603_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X139 a_1393_1862# a_1293_1765# a_1235_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X140 a_n503_n2934# a_n603_n3031# a_n661_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X141 a_n661_n1626# a_n761_n1723# a_n819_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X142 a_n1293_1862# a_n1393_1765# a_n1451_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X143 a_n503_n1190# a_n603_n1287# a_n661_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X144 a_n1451_990# a_n1551_893# a_n1609_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X145 a_445_1426# a_345_1329# a_287_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X146 a_287_n2934# a_187_n3031# a_129_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X147 a_761_n2062# a_661_n2159# a_603_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X148 a_287_n1190# a_187_n1287# a_129_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X149 a_129_2734# a_29_2637# a_n29_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X150 a_n345_n318# a_n445_n415# a_n503_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X151 a_n1451_1426# a_n1551_1329# a_n1609_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X152 a_1551_1426# a_1451_1329# a_1393_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X153 a_n661_554# a_n761_457# a_n819_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X154 a_n661_n2934# a_n761_n3031# a_n819_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X155 a_n345_2298# a_n445_2201# a_n503_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X156 a_n503_118# a_n603_21# a_n661_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X157 a_n1135_n1626# a_n1235_n1723# a_n1293_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X158 a_n661_n1190# a_n761_n1287# a_n819_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X159 a_129_554# a_29_457# a_n29_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X160 a_n503_n2498# a_n603_n2595# a_n661_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X161 a_445_2734# a_345_2637# a_287_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X162 a_n977_990# a_n1077_893# a_n1135_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X163 a_287_n754# a_187_n851# a_129_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X164 a_129_n318# a_29_n415# a_n29_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X165 a_287_n2498# a_187_n2595# a_129_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X166 a_1551_2734# a_1451_2637# a_1393_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X167 a_n1451_2734# a_n1551_2637# a_n1609_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X168 a_129_2298# a_29_2201# a_n29_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X169 a_n187_554# a_n287_457# a_n345_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X170 a_n1293_n754# a_n1393_n851# a_n1451_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X171 a_1393_n754# a_1293_n851# a_1235_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X172 a_n1293_n1626# a_n1393_n1723# a_n1451_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X173 a_n29_118# a_n129_21# a_n187_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X174 a_n1135_n1190# a_n1235_n1287# a_n1293_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X175 a_n1135_n2934# a_n1235_n3031# a_n1293_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X176 a_n661_n2498# a_n761_n2595# a_n819_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X177 a_n345_1862# a_n445_1765# a_n503_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X178 a_445_n318# a_345_n415# a_287_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X179 a_1551_n1626# a_1451_n1723# a_1393_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X180 a_n29_n1626# a_n129_n1723# a_n187_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X181 a_445_2298# a_345_2201# a_287_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X182 a_n977_1426# a_n1077_1329# a_n1135_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X183 a_n1135_990# a_n1235_893# a_n1293_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X184 a_1551_n318# a_1451_n415# a_1393_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X185 a_n1451_n318# a_n1551_n415# a_n1609_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X186 a_1551_2298# a_1451_2201# a_1393_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X187 a_1077_1426# a_977_1329# a_919_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X188 a_n819_554# a_n919_457# a_n977_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X189 a_1393_118# a_1293_21# a_1235_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X190 a_n1293_n2934# a_n1393_n3031# a_n1451_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X191 a_n1451_2298# a_n1551_2201# a_n1609_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X192 a_n503_1426# a_n603_1329# a_n661_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X193 a_n345_554# a_n445_457# a_n503_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X194 a_n1293_n1190# a_n1393_n1287# a_n1451_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X195 a_n1135_n2498# a_n1235_n2595# a_n1293_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X196 a_129_1862# a_29_1765# a_n29_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X197 a_n29_n2934# a_n129_n3031# a_n187_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X198 a_n187_n1626# a_n287_n1723# a_n345_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X199 a_n977_2734# a_n1077_2637# a_n1135_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X200 a_1551_n2934# a_1451_n3031# a_1393_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X201 a_n503_n2062# a_n603_n2159# a_n661_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X202 a_n29_n1190# a_n129_n1287# a_n187_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X203 a_1551_n1190# a_1451_n1287# a_1393_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X204 a_1077_118# a_977_21# a_919_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X205 a_1077_2734# a_977_2637# a_919_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X206 a_445_1862# a_345_1765# a_287_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X207 a_287_n2062# a_187_n2159# a_129_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X208 a_n503_2734# a_n603_2637# a_n661_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X209 a_n345_n754# a_n445_n851# a_n503_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X210 a_n1293_n2498# a_n1393_n2595# a_n1451_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X211 a_n1451_1862# a_n1551_1765# a_n1609_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X212 a_1551_1862# a_1451_1765# a_1393_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X213 a_n661_990# a_n761_893# a_n819_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X214 a_1551_118# a_1451_21# a_1393_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X215 a_n977_n318# a_n1077_n415# a_n1135_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X216 a_n187_n2934# a_n287_n3031# a_n345_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X217 a_n661_n2062# a_n761_n2159# a_n819_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X218 a_n503_554# a_n603_457# a_n661_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X219 a_1551_n2498# a_1451_n2595# a_1393_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X220 a_n29_n2498# a_n129_n2595# a_n187_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X221 a_n187_n1190# a_n287_n1287# a_n345_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X222 a_n977_2298# a_n1077_2201# a_n1135_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X223 a_n29_1426# a_n129_1329# a_n187_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X224 a_603_1426# a_503_1329# a_445_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X225 a_129_990# a_29_893# a_n29_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X226 a_1077_n318# a_977_n415# a_919_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X227 a_n503_n318# a_n603_n415# a_n661_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X228 a_1077_2298# a_977_2201# a_919_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X229 a_129_n754# a_29_n851# a_n29_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X230 a_n503_2298# a_n603_2201# a_n661_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X231 a_761_118# a_661_21# a_603_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X232 a_n187_990# a_n287_893# a_n345_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X233 a_n187_n2498# a_n287_n2595# a_n345_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X234 a_n1135_n2062# a_n1235_n2159# a_n1293_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X235 a_n29_554# a_n129_457# a_n187_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X236 a_129_n1626# a_29_n1723# a_n29_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X237 a_n29_2734# a_n129_2637# a_n187_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X238 a_603_2734# a_503_2637# a_445_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X239 a_445_n754# a_345_n851# a_287_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X240 a_n977_1862# a_n1077_1765# a_n1135_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X241 a_1551_n754# a_1451_n851# a_1393_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X242 a_287_118# a_187_21# a_129_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X243 a_n1451_n754# a_n1551_n851# a_n1609_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X244 a_1077_1862# a_977_1765# a_919_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X245 a_n819_990# a_n919_893# a_n977_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X246 a_1393_554# a_1293_457# a_1235_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X247 a_n1293_n2062# a_n1393_n2159# a_n1451_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X248 a_n503_1862# a_n603_1765# a_n661_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X249 a_1235_118# a_1135_21# a_1077_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X250 a_n29_n318# a_n129_n415# a_n187_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X251 a_603_n318# a_503_n415# a_445_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X252 a_129_n2934# a_29_n3031# a_n29_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X253 a_603_2298# a_503_2201# a_445_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X254 a_n1135_1426# a_n1235_1329# a_n1293_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X255 a_1235_1426# a_1135_1329# a_1077_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X256 a_n345_990# a_n445_893# a_n503_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X257 a_1551_n2062# a_1451_n2159# a_1393_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X258 a_n29_n2062# a_n129_n2159# a_n187_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X259 a_129_n1190# a_29_n1287# a_n29_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X260 a_n29_2298# a_n129_2201# a_n187_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X261 a_445_n1626# a_345_n1723# a_287_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X262 a_1077_554# a_977_457# a_919_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X263 a_919_118# a_819_21# a_761_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X264 a_1235_2734# a_1135_2637# a_1077_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X265 a_445_118# a_345_21# a_287_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X266 a_129_n2498# a_29_n2595# a_n29_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X267 a_n187_n2062# a_n287_n2159# a_n345_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X268 a_n1135_2734# a_n1235_2637# a_n1293_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X269 a_1551_554# a_1451_457# a_1393_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X270 a_n977_n754# a_n1077_n851# a_n1135_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X271 a_n503_990# a_n603_893# a_n661_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X272 a_445_n2934# a_345_n3031# a_287_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X273 a_n29_1862# a_n129_1765# a_n187_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X274 a_603_1862# a_503_1765# a_445_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X275 a_445_n1190# a_345_n1287# a_287_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X276 a_1077_n754# a_977_n851# a_919_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X277 a_n503_n754# a_n603_n851# a_n661_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X278 a_919_n1626# a_819_n1723# a_761_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X279 a_1235_n318# a_1135_n415# a_1077_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQFY a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQ24 a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt follower_amp vdd out ena in vsub vss
XXM12 m1_651_3930# m1_651_3930# out m1_651_3930# vdd out vdd m1_651_3930# vdd out
+ vdd out out m1_651_3930# out vdd m1_651_3930# m1_651_3930# vdd vdd out m1_651_3930#
+ m1_651_3930# out m1_651_3930# m1_651_3930# out vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ out m1_651_3930# m1_651_3930# vdd vdd vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ m1_651_3930# out sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW
XXM13 m1_2399_1244# vss nbias ena sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM24 pbias vss vss nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM25 pbias vdd pbias vcomp vdd vdd pbias pbias sky130_fd_pr__pfet_g5v0d10v5_KLJMY6
XXM27 vcomp m2_526_2596# vdd vcomp out in out m1_811_2614# in vcomp sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXM29 m1_811_2614# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXR1 m1_3337_606# vdd m1_604_772# m1_604_772# m1_2399_1244# m1_3337_606# vss sky130_fd_pr__res_xhigh_po_0p35_HLA228
XXM1 vss m2_1742_2323# m1_505_3709# m2_1930_2454# out in sky130_fd_pr__nfet_g5v0d10v5_FJGQFC
XXM5 vdd m1_505_3709# vdd vdd m2_1930_2454# m2_1930_2454# m2_1930_2454# m2_1930_2454#
+ m2_1930_2454# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXXD1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__1
XXM6 vdd m1_651_3930# vdd vdd m2_3105_2460# m2_3105_2460# m2_3105_2460# m2_3105_2460#
+ m2_3105_2460# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXXD2 vss in sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__1
XXM7 vss vss m2_2845_2323# m2_2845_2323# nbias nbias sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y
XXM8 vss vss m2_1742_2323# nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM9 m2_2845_2323# m2_3105_2460# in vss m1_651_3930# out sky130_fd_pr__nfet_05v0_nvt_BH6ZTK
XXM30 m2_526_2596# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM20 out vdd m1_505_3709# out vdd out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd m1_505_3709# out vdd m1_505_3709# out m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd out m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ vdd out vdd m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# out out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# out out out m1_505_3709# m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd out vdd m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out out m1_505_3709# vdd out
+ out out m1_505_3709# vdd vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# out m1_505_3709# vdd m1_505_3709# out
+ m1_505_3709# m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# out vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd out vdd
+ vdd m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# out m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# out out vdd out m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# out out vdd vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709# vdd out vdd out
+ out m1_505_3709# vdd vdd out out out m1_505_3709# m1_505_3709# m1_505_3709# out
+ out vdd out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd vdd out vdd m1_505_3709# vdd
+ out out m1_505_3709# out m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out vdd m1_505_3709#
+ m1_505_3709# vdd out vdd out m1_505_3709# out m1_505_3709# out m1_505_3709# out
+ m1_505_3709# vdd m1_505_3709# out m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd vdd m1_505_3709# m1_505_3709# out vdd vdd vdd
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# out vdd out out m1_505_3709# out out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd out vdd out m1_505_3709# vdd out m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out vdd out vdd
+ out m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# out m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# vdd out out m1_505_3709# vdd vdd out out vdd m1_505_3709#
+ out m1_505_3709# vdd out m1_505_3709# m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out out vdd m1_505_3709#
+ vdd out m1_505_3709# out vdd out m1_505_3709# vdd out out vdd out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# out vdd vdd out vdd out out m1_505_3709# vdd m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# vdd out
+ m1_505_3709# m1_505_3709# out sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ
XXM10 nbias vss nbias vss nbias vss vss nbias nbias nbias sky130_fd_pr__nfet_g5v0d10v5_H7BQFY
XXM22 m2_526_2596# vss out vss out vss vss m2_526_2596# m2_526_2596# m2_526_2596#
+ sky130_fd_pr__nfet_g5v0d10v5_H7BQ24
.ends

.subckt dac_3v_column b4b dum1_out b0_uq12 b0_uq1 b2b_uq0 dac_3v_cell_top_0/m4_97_801#
+ b0_uq11 b0_uq10 b2b_uq2 b3b b4 b0b_uq13 b2b_uq1 b0_uq6 dac_3v_cell_0[2]/w_316_892#
+ dum0_in dac_3v_cell_0[1]/w_316_892# b0b_uq11 b0 dac_3v_cell_top_0/m4_97_1059# b1
+ b0b_uq10 b1_uq6 dac_3v_cell_0[6]/w_316_892# b0b_uq12 b1_uq1 b1_uq2 b1_uq0 b3 b0_uq3
+ b0b_uq2 b1_uq3 b0b_uq1 b0_uq14 dac_3v_cell_0[5]/w_316_892# b0b_uq14 b0b_uq7 b0b_uq0
+ b0_uq2 b0b_uq6 out_5 b0b_uq9 out_4 dac_3v_cell_top_0/m1_290_591# b0b_uq8 b1b_uq6
+ b0_uq13 b3_uq0 b3b_uq0 b1b_uq5 dac_3v_cell_0[4]/w_316_892# b2_uq1 res0_in b2 m2_801_196#
+ b1b_uq4 b0_uq5 b0_uq0 b2_uq0 b1b_uq3 b0_uq4 b1b_uq2 b1_uq5 b2_uq2 m2_791_1314# b1_uq4
+ b1b_uq0 b0b_uq5 m2_791_14877# dac_3v_cell_0[7]/w_316_892# b0_uq9 b0b b1b_uq1 res1_out
+ dac_3v_cell_top_0/m1_290_1114# b0_uq8 dac_3v_cell_0[3]/w_316_892# b1b b0b_uq4 b0b_uq3
+ b0_uq7 m2_801_13759# b2b VSUBS
Xdac_3v_cell_0[0] m2_791_1314# m2_801_196# m2_328_1119# m2_328_1119# res1_out m2_791_1314#
+ VSUBS m2_449_485# m2_328_1119# dum1_out m2_801_196# m2_449_485# VSUBS m2_449_485#
+ VSUBS m2_791_1314# m2_801_196# VSUBS res0_in dum0_in VSUBS dac_3v_cell
Xdac_3v_cell_0[1] b0b m2_791_1314# out0_0_0 out0_1_0 dac_3v_cell_0[1]/m1_824_799#
+ b1b_uq0 VSUBS out0_0_0 out1_0_3 res1_out b0_uq0 out_3 b4b out_4 b0 dac_3v_cell_0[1]/w_316_892#
+ b4 b1_uq0 dac_3v_cell_0[2]/m1_155_n223# res0_in b0b_uq0 dac_3v_cell
Xdac_3v_cell_0[2] b0_uq2 dac_3v_cell_0[1]/w_316_892# out0_2 out0_1_0 dac_3v_cell_0[2]/m1_824_799#
+ b2b_uq0 VSUBS out0_0_0 out1_0_3 dac_3v_cell_0[1]/m1_824_799# b0b_uq1 out1_1_1 b1b
+ out1_0_3 b0b_uq2 dac_3v_cell_0[2]/w_316_892# b1 b2_uq0 dac_3v_cell_0[3]/m1_155_n223#
+ dac_3v_cell_0[2]/m1_155_n223# b0_uq1 dac_3v_cell
Xdac_3v_cell_0[3] b0b_uq4 dac_3v_cell_0[2]/w_316_892# out0_0_1 out0_1_0 dac_3v_cell_0[3]/m1_824_799#
+ b1_uq1 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[2]/m1_824_799# b0_uq3 out1_1_1 b2b
+ out1_2 b0_uq4 dac_3v_cell_0[3]/w_316_892# b2 b1b_uq1 dac_3v_cell_0[4]/m1_155_n223#
+ dac_3v_cell_0[3]/m1_155_n223# b0b_uq3 dac_3v_cell
Xdac_3v_cell_0[4] b0_uq6 dac_3v_cell_0[3]/w_316_892# out_3 out0_2 dac_3v_cell_0[4]/m1_824_799#
+ b3b_uq0 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[3]/m1_824_799# b0b_uq5 out1_1_1 b1_uq2
+ out1_0_2 b0b_uq6 dac_3v_cell_0[4]/w_316_892# b1b_uq2 b3_uq0 dac_3v_cell_0[5]/m1_155_n223#
+ dac_3v_cell_0[4]/m1_155_n223# b0_uq5 dac_3v_cell
Xdac_3v_cell_0[5] b0b_uq8 dac_3v_cell_0[4]/w_316_892# out0_0_2 out0_1_1 dac_3v_cell_0[5]/m1_824_799#
+ b1b_uq3 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[4]/m1_824_799# b0_uq7 out1_2 b3b out_3
+ b0_uq8 dac_3v_cell_0[5]/w_316_892# b3 b1_uq3 dac_3v_cell_0[6]/m1_155_n223# dac_3v_cell_0[5]/m1_155_n223#
+ b0b_uq7 dac_3v_cell
Xdac_3v_cell_0[6] b0_uq10 dac_3v_cell_0[5]/w_316_892# out0_2 out0_1_1 dac_3v_cell_0[6]/m1_824_799#
+ b2_uq1 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[5]/m1_824_799# b0b_uq9 out1_1_0 b1b_uq4
+ out1_0_1 b0b_uq10 dac_3v_cell_0[6]/w_316_892# b1_uq4 b2b_uq1 dac_3v_cell_0[7]/m1_155_n223#
+ dac_3v_cell_0[6]/m1_155_n223# b0_uq9 dac_3v_cell
Xdac_3v_cell_0[7] b0b_uq12 dac_3v_cell_0[6]/w_316_892# out0_0_3 out0_1_1 dac_3v_cell_0[7]/m1_824_799#
+ b1_uq5 VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[6]/m1_824_799# b0_uq11 out1_1_0 b2_uq2
+ out1_2 b0_uq12 dac_3v_cell_0[7]/w_316_892# b2b_uq2 b1b_uq5 dac_3v_cell_top_0/m1_155_n223#
+ dac_3v_cell_0[7]/m1_155_n223# b0b_uq11 dac_3v_cell
Xdac_3v_cell_1 m2_791_14877# m2_801_13759# m2_330_14682# m2_330_14682# dum0_out m2_791_14877#
+ VSUBS m2_449_14048# m2_330_14682# res1_in m2_801_13759# m2_449_14048# VSUBS m2_449_14048#
+ VSUBS m2_791_14877# m2_801_13759# VSUBS dum0_out res1_in VSUBS dac_3v_cell
Xdac_3v_cell_top_0 b0_uq14 dac_3v_cell_0[7]/w_316_892# out_4 out_5 res1_in m2_801_13759#
+ dac_3v_cell_top_0/m1_290_1114# VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[7]/m1_824_799#
+ b0b_uq13 dac_3v_cell_top_0/m4_97_801# out1_1_0 dac_3v_cell_top_0/m4_97_1059# b1_uq6
+ out1_0_0 b0b_uq14 b1b_uq6 dac_3v_cell_top_0/m1_290_591# dac_3v_cell_top_0/m1_155_n223#
+ b0_uq13 dac_3v_cell_top
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_4AXGXB a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt rdac_level_shifter dvdd bitb_out bit_out bit_in avdd agnd
Xsky130_fd_sc_hvl__inv_8_1 bitb_out agnd agnd avdd avdd bit_out sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 bit_in dvdd agnd avdd avdd sky130_fd_sc_hvl__inv_2_0/A
+ avdd agnd agnd sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_4AXGXB_0 agnd bit_in sky130_fd_pr__diode_pw2nd_05v5_4AXGXB
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A agnd agnd avdd avdd bitb_out
+ sky130_fd_sc_hvl__inv_8
.ends

.subckt level_shifter_array rdac_level_shifter_0[2]/bit_out rdac_level_shifter_0[6]/bitb_out
+ rdac_level_shifter_0[2]/bitb_out rdac_level_shifter_0[3]/bit_in rdac_level_shifter_0[7]/bit_in
+ rdac_level_shifter_0[6]/bit_out rdac_level_shifter_0[3]/bit_out rdac_level_shifter_0[7]/dvdd
+ rdac_level_shifter_0[0]/bit_in rdac_level_shifter_0[3]/bitb_out rdac_level_shifter_0[0]/bit_out
+ rdac_level_shifter_0[4]/bit_in rdac_level_shifter_0[7]/bit_out rdac_level_shifter_0[4]/bit_out
+ rdac_level_shifter_0[4]/bitb_out rdac_level_shifter_0[1]/bit_in rdac_level_shifter_0[0]/bitb_out
+ rdac_level_shifter_0[5]/bit_in rdac_level_shifter_0[1]/bit_out rdac_level_shifter_0[7]/bitb_out
+ rdac_level_shifter_0[5]/bitb_out rdac_level_shifter_0[5]/bit_out rdac_level_shifter_0[2]/bit_in
+ rdac_level_shifter_0[1]/bitb_out VSUBS rdac_level_shifter_0[6]/bit_in rdac_level_shifter_0[7]/avdd
Xrdac_level_shifter_0[0] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[0]/bitb_out
+ rdac_level_shifter_0[0]/bit_out rdac_level_shifter_0[0]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[1] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[1]/bitb_out
+ rdac_level_shifter_0[1]/bit_out rdac_level_shifter_0[1]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[2] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[2]/bitb_out
+ rdac_level_shifter_0[2]/bit_out rdac_level_shifter_0[2]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[3] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[3]/bitb_out
+ rdac_level_shifter_0[3]/bit_out rdac_level_shifter_0[3]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[4] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[4]/bitb_out
+ rdac_level_shifter_0[4]/bit_out rdac_level_shifter_0[4]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[5] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[5]/bitb_out
+ rdac_level_shifter_0[5]/bit_out rdac_level_shifter_0[5]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[6] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[6]/bitb_out
+ rdac_level_shifter_0[6]/bit_out rdac_level_shifter_0[6]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[7] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[7]/bitb_out
+ rdac_level_shifter_0[7]/bit_out rdac_level_shifter_0[7]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
.ends

.subckt dac_3v_cell_dummy m4_99_18# w_318_n275# m4_99_276# m4_99_801# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m4_99_930# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m4_99_405# m4_99_1059#
+ m4_99_672# w_316_892# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300# m4_99_147#
+ m1_155_n223# m1_824_799#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_387_847# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_545_212# m1_545_212# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt dac_3v_column_dummy m1_988_1608# dac_3v_cell_dummy_0[6]/m4_99_147# dac_3v_cell_dummy_0[0]/w_318_n275#
+ dac_3v_cell_dummy_0[7]/m4_99_147# dac_3v_cell_dummy_0[6]/m4_99_18# dac_3v_cell_dummy_0[8]/m4_99_147#
+ dac_3v_cell_dummy_0[9]/m4_99_147# dac_3v_cell_dummy_0[7]/m4_99_18# dac_3v_cell_dummy_0[0]/m4_99_276#
+ dac_3v_cell_dummy_0[0]/m4_99_801# dac_3v_cell_dummy_0[1]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_1059#
+ dac_3v_cell_dummy_0[2]/m4_99_1059# dac_3v_cell_dummy_0[1]/m4_99_801# dac_3v_cell_dummy_0[2]/m4_99_276#
+ dac_3v_cell_dummy_0[2]/m4_99_801# dac_3v_cell_dummy_0[3]/m4_99_276# dac_3v_cell_dummy_0[3]/m4_99_801#
+ dac_3v_cell_dummy_0[4]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_18# dac_3v_cell_dummy_0[4]/m4_99_801#
+ dac_3v_cell_dummy_0[5]/m4_99_276# dac_3v_cell_dummy_0[5]/m4_99_801# dac_3v_cell_dummy_0[6]/m4_99_276#
+ dac_3v_cell_dummy_0[6]/m4_99_801# dac_3v_cell_dummy_0[7]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_801#
+ dac_3v_cell_dummy_0[9]/m4_99_18# dac_3v_cell_dummy_0[8]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_801#
+ dac_3v_cell_dummy_0[9]/m4_99_276# dac_3v_cell_dummy_0[9]/m4_99_801# dac_3v_cell_dummy_0[6]/m4_99_1059#
+ dac_3v_cell_dummy_0[1]/m4_99_1059# dac_3v_cell_dummy_0[0]/m4_99_930# dac_3v_cell_dummy_0[1]/m4_99_930#
+ dac_3v_cell_dummy_0[2]/m4_99_930# dac_3v_cell_dummy_0[3]/m4_99_930# dac_3v_cell_dummy_0[0]/m4_99_18#
+ dac_3v_cell_dummy_0[4]/m4_99_930# dac_3v_cell_dummy_0[5]/m4_99_930# dac_3v_cell_dummy_0[6]/m4_99_930#
+ VSUBS dac_3v_cell_dummy_0[5]/m4_99_1059# dac_3v_cell_dummy_0[7]/m4_99_930# dac_3v_cell_dummy_0[1]/m4_99_18#
+ dac_3v_cell_dummy_0[0]/m4_99_1059# dac_3v_cell_dummy_0[8]/m4_99_930# dac_3v_cell_dummy_0[9]/m4_99_930#
+ dac_3v_cell_dummy_0[0]/m4_99_405# dac_3v_cell_dummy_0[1]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_405#
+ dac_3v_cell_dummy_0[0]/m4_99_672# dac_3v_cell_dummy_0[2]/m4_99_18# dac_3v_cell_dummy_0[3]/m4_99_405#
+ m1_938_45# dac_3v_cell_dummy_0[1]/m4_99_672# dac_3v_cell_dummy_0[4]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_672#
+ dac_3v_cell_dummy_0[1]/w_316_892# dac_3v_cell_dummy_0[5]/m4_99_405# dac_3v_cell_dummy_0[3]/m4_99_672#
+ dac_3v_cell_dummy_0[2]/w_316_892# dac_3v_cell_dummy_0[4]/m4_99_672# dac_3v_cell_dummy_0[6]/m4_99_405#
+ dac_3v_cell_dummy_0[9]/m4_99_1059# dac_3v_cell_dummy_0[3]/m4_99_18# dac_3v_cell_dummy_0[4]/m4_99_1059#
+ dac_3v_cell_dummy_0[3]/w_316_892# dac_3v_cell_dummy_0[5]/m4_99_672# dac_3v_cell_dummy_0[7]/m4_99_405#
+ dac_3v_cell_dummy_0[8]/m4_99_405# dac_3v_cell_dummy_0[6]/m4_99_672# dac_3v_cell_dummy_0[4]/w_316_892#
+ dac_3v_cell_dummy_0[0]/w_316_892# dac_3v_cell_dummy_0[7]/m4_99_672# dac_3v_cell_dummy_0[9]/m4_99_405#
+ dac_3v_cell_dummy_0[5]/w_316_892# dac_3v_cell_dummy_0[6]/w_316_892# dac_3v_cell_dummy_0[8]/m4_99_672#
+ dac_3v_cell_dummy_0[4]/m4_99_18# dac_3v_cell_dummy_0[7]/w_316_892# dac_3v_cell_dummy_0[0]/m4_99_147#
+ dac_3v_cell_dummy_0[9]/m4_99_672# dac_3v_cell_dummy_0[8]/w_316_892# dac_3v_cell_dummy_0[1]/m4_99_147#
+ m1_n18_1607# dac_3v_cell_dummy_0[9]/w_316_892# dac_3v_cell_dummy_0[2]/m4_99_147#
+ dac_3v_cell_dummy_0[3]/m4_99_147# dac_3v_cell_dummy_0[5]/m4_99_18# m1_n18_45# dac_3v_cell_dummy_0[8]/m4_99_1059#
+ dac_3v_cell_dummy_0[4]/m4_99_147# dac_3v_cell_dummy_0[3]/m4_99_1059# dac_3v_cell_dummy_0[5]/m4_99_147#
Xdac_3v_cell_dummy_0[0] dac_3v_cell_dummy_0[0]/m4_99_18# dac_3v_cell_dummy_0[0]/w_318_n275#
+ dac_3v_cell_dummy_0[0]/m4_99_276# dac_3v_cell_dummy_0[0]/m4_99_801# VSUBS dac_3v_cell_dummy_0[0]/m4_99_930#
+ m1_938_45# dac_3v_cell_dummy_0[0]/m4_99_405# dac_3v_cell_dummy_0[0]/m4_99_1059#
+ dac_3v_cell_dummy_0[0]/m4_99_672# dac_3v_cell_dummy_0[0]/w_316_892# m1_n18_1607#
+ dac_3v_cell_dummy_0[0]/m4_99_147# m1_n18_45# m1_988_1608# dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[1] dac_3v_cell_dummy_0[1]/m4_99_18# dac_3v_cell_dummy_0[0]/w_316_892#
+ dac_3v_cell_dummy_0[1]/m4_99_276# dac_3v_cell_dummy_0[1]/m4_99_801# VSUBS dac_3v_cell_dummy_0[1]/m4_99_930#
+ m1_988_1608# dac_3v_cell_dummy_0[1]/m4_99_405# dac_3v_cell_dummy_0[1]/m4_99_1059#
+ dac_3v_cell_dummy_0[1]/m4_99_672# dac_3v_cell_dummy_0[1]/w_316_892# dac_3v_cell_dummy_0[2]/m1_155_n223#
+ dac_3v_cell_dummy_0[1]/m4_99_147# m1_n18_1607# dac_3v_cell_dummy_0[1]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[2] dac_3v_cell_dummy_0[2]/m4_99_18# dac_3v_cell_dummy_0[1]/w_316_892#
+ dac_3v_cell_dummy_0[2]/m4_99_276# dac_3v_cell_dummy_0[2]/m4_99_801# VSUBS dac_3v_cell_dummy_0[2]/m4_99_930#
+ dac_3v_cell_dummy_0[1]/m1_824_799# dac_3v_cell_dummy_0[2]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_1059#
+ dac_3v_cell_dummy_0[2]/m4_99_672# dac_3v_cell_dummy_0[2]/w_316_892# dac_3v_cell_dummy_0[3]/m1_155_n223#
+ dac_3v_cell_dummy_0[2]/m4_99_147# dac_3v_cell_dummy_0[2]/m1_155_n223# dac_3v_cell_dummy_0[2]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[3] dac_3v_cell_dummy_0[3]/m4_99_18# dac_3v_cell_dummy_0[2]/w_316_892#
+ dac_3v_cell_dummy_0[3]/m4_99_276# dac_3v_cell_dummy_0[3]/m4_99_801# VSUBS dac_3v_cell_dummy_0[3]/m4_99_930#
+ dac_3v_cell_dummy_0[2]/m1_824_799# dac_3v_cell_dummy_0[3]/m4_99_405# dac_3v_cell_dummy_0[3]/m4_99_1059#
+ dac_3v_cell_dummy_0[3]/m4_99_672# dac_3v_cell_dummy_0[3]/w_316_892# dac_3v_cell_dummy_0[4]/m1_155_n223#
+ dac_3v_cell_dummy_0[3]/m4_99_147# dac_3v_cell_dummy_0[3]/m1_155_n223# dac_3v_cell_dummy_0[3]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[4] dac_3v_cell_dummy_0[4]/m4_99_18# dac_3v_cell_dummy_0[3]/w_316_892#
+ dac_3v_cell_dummy_0[4]/m4_99_276# dac_3v_cell_dummy_0[4]/m4_99_801# VSUBS dac_3v_cell_dummy_0[4]/m4_99_930#
+ dac_3v_cell_dummy_0[3]/m1_824_799# dac_3v_cell_dummy_0[4]/m4_99_405# dac_3v_cell_dummy_0[4]/m4_99_1059#
+ dac_3v_cell_dummy_0[4]/m4_99_672# dac_3v_cell_dummy_0[4]/w_316_892# dac_3v_cell_dummy_0[5]/m1_155_n223#
+ dac_3v_cell_dummy_0[4]/m4_99_147# dac_3v_cell_dummy_0[4]/m1_155_n223# dac_3v_cell_dummy_0[4]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[5] dac_3v_cell_dummy_0[5]/m4_99_18# dac_3v_cell_dummy_0[4]/w_316_892#
+ dac_3v_cell_dummy_0[5]/m4_99_276# dac_3v_cell_dummy_0[5]/m4_99_801# VSUBS dac_3v_cell_dummy_0[5]/m4_99_930#
+ dac_3v_cell_dummy_0[4]/m1_824_799# dac_3v_cell_dummy_0[5]/m4_99_405# dac_3v_cell_dummy_0[5]/m4_99_1059#
+ dac_3v_cell_dummy_0[5]/m4_99_672# dac_3v_cell_dummy_0[5]/w_316_892# dac_3v_cell_dummy_0[6]/m1_155_n223#
+ dac_3v_cell_dummy_0[5]/m4_99_147# dac_3v_cell_dummy_0[5]/m1_155_n223# dac_3v_cell_dummy_0[5]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[6] dac_3v_cell_dummy_0[6]/m4_99_18# dac_3v_cell_dummy_0[5]/w_316_892#
+ dac_3v_cell_dummy_0[6]/m4_99_276# dac_3v_cell_dummy_0[6]/m4_99_801# VSUBS dac_3v_cell_dummy_0[6]/m4_99_930#
+ dac_3v_cell_dummy_0[5]/m1_824_799# dac_3v_cell_dummy_0[6]/m4_99_405# dac_3v_cell_dummy_0[6]/m4_99_1059#
+ dac_3v_cell_dummy_0[6]/m4_99_672# dac_3v_cell_dummy_0[6]/w_316_892# dac_3v_cell_dummy_0[7]/m1_155_n223#
+ dac_3v_cell_dummy_0[6]/m4_99_147# dac_3v_cell_dummy_0[6]/m1_155_n223# dac_3v_cell_dummy_0[6]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[7] dac_3v_cell_dummy_0[7]/m4_99_18# dac_3v_cell_dummy_0[6]/w_316_892#
+ dac_3v_cell_dummy_0[7]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_801# VSUBS dac_3v_cell_dummy_0[7]/m4_99_930#
+ dac_3v_cell_dummy_0[6]/m1_824_799# dac_3v_cell_dummy_0[7]/m4_99_405# dac_3v_cell_dummy_0[7]/m4_99_1059#
+ dac_3v_cell_dummy_0[7]/m4_99_672# dac_3v_cell_dummy_0[7]/w_316_892# dac_3v_cell_dummy_0[8]/m1_155_n223#
+ dac_3v_cell_dummy_0[7]/m4_99_147# dac_3v_cell_dummy_0[7]/m1_155_n223# dac_3v_cell_dummy_0[7]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[8] dac_3v_cell_dummy_0[8]/m4_99_18# dac_3v_cell_dummy_0[7]/w_316_892#
+ dac_3v_cell_dummy_0[8]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_801# VSUBS dac_3v_cell_dummy_0[8]/m4_99_930#
+ dac_3v_cell_dummy_0[7]/m1_824_799# dac_3v_cell_dummy_0[8]/m4_99_405# dac_3v_cell_dummy_0[8]/m4_99_1059#
+ dac_3v_cell_dummy_0[8]/m4_99_672# dac_3v_cell_dummy_0[8]/w_316_892# m1_36_13186#
+ dac_3v_cell_dummy_0[8]/m4_99_147# dac_3v_cell_dummy_0[8]/m1_155_n223# m1_36_13186#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[9] dac_3v_cell_dummy_0[9]/m4_99_18# dac_3v_cell_dummy_0[8]/w_316_892#
+ dac_3v_cell_dummy_0[9]/m4_99_276# dac_3v_cell_dummy_0[9]/m4_99_801# VSUBS dac_3v_cell_dummy_0[9]/m4_99_930#
+ m1_36_13186# dac_3v_cell_dummy_0[9]/m4_99_405# dac_3v_cell_dummy_0[9]/m4_99_1059#
+ dac_3v_cell_dummy_0[9]/m4_99_672# dac_3v_cell_dummy_0[9]/w_316_892# m1_28_15111#
+ dac_3v_cell_dummy_0[9]/m4_99_147# m1_36_13186# m1_28_15111# dac_3v_cell_dummy
.ends

.subckt sky130_ef_ip__rdac3v_8bit b0 b1 b2 b3 b4 b5 b6 b7 out vdd ena dvdd Vhigh Vlow
+ vss dvss
Xdac_3v_column_odd_0 b6b dac_3v_column_0/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_1/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_0/dum1_out b0a b1a dac_3v_column_1/res0_in b0b b2b b2a dac_3v_column_0/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_1/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_1 b7b dac_3v_column_1/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b7a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a out_unbuf b1b b1b b3a vdd vdd dac_3v_column_1/dum1_out
+ b0a b1a dac_3v_column_2/res0_in b0b b2b b2a dac_3v_column_1/out_4 b1a vdd b2b b3b
+ vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_2/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_2 b6a dac_3v_column_2/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_3/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_2/dum1_out b0a b1a dac_3v_column_3/res0_in b0b b2b b2a dac_3v_column_2/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_3/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_3 vdd dac_3v_column_3/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a vss b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_odd_3/in_5 b1b b1b b3a vdd
+ vdd dac_3v_column_3/dum1_out b0a b1a dac_3v_column_4/res0_in b0b b2b b2a dac_3v_column_3/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_3/in_5
+ b0a dac_3v_column_4/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_4 b6b dac_3v_column_4/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_5/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_4/dum1_out b0a b1a dac_3v_column_5/res0_in b0b b2b b2a dac_3v_column_4/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_5/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xfollower_amp_0 vdd out ena out_unbuf dvss vss follower_amp
Xdac_3v_column_odd_5 b7a dac_3v_column_5/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b7b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a out_unbuf b1b b1b b3a vdd vdd dac_3v_column_5/dum1_out
+ b0a b1a dac_3v_column_6/res0_in b0b b2b b2a dac_3v_column_5/out_4 b1a vdd b2b b3b
+ vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_6/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_6 b6a dac_3v_column_6/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_7/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_6/dum1_out b0a b1a dac_3v_column_7/res0_in b0b b2b b2a dac_3v_column_6/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_7/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_7 vdd dac_3v_column_7/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a vss b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_odd_7/in_5 b1b b1b b3a vdd
+ vdd dac_3v_column_7/dum1_out b0a b1a Vlow b0b b2b b2a dac_3v_column_7/out_4 b1a
+ vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_7/in_5
+ b0a dac_3v_column_odd_7/dum_out1 b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_0 b4b dac_3v_column_0/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_0/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_1/out_5 b0a
+ dac_3v_column_0/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b Vhigh b2b vdd b1a b0b
+ b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a dac_3v_column_0/res1_out
+ b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_1 b4b dac_3v_column_1/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_1/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_1/out_5 b0a
+ dac_3v_column_1/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_1/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_1/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_2 b4b dac_3v_column_2/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_2/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_3/out_5 b0a
+ dac_3v_column_2/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_2/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_2/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_3 b4b dac_3v_column_3/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_3/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_3/out_5 b0a
+ dac_3v_column_3/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_3/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_3/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_4 b4b dac_3v_column_4/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_4/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_5/out_5 b0a
+ dac_3v_column_4/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_4/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_4/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_5 b4b dac_3v_column_5/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_5/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_5/out_5 b0a
+ dac_3v_column_5/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_5/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_5/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_6 b4b dac_3v_column_6/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_6/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_7/out_5 b0a
+ dac_3v_column_6/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_6/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_6/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_7 b4b dac_3v_column_7/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_7/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_7/out_5 b0a
+ dac_3v_column_7/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_7/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_7/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xlevel_shifter_array_0 b2b b6b b2a b3 b7 b6a b3b dvdd b0 b3a b0a b4 b7a b4b b4a b1
+ b0b b5 b1b b7b b5a b5b b2 b1a dvss b6 vdd level_shifter_array
Xdac_3v_column_dummy_0 Vhigh b0a vdd b0b b1b b0a vdd b2a vss vss b4b b1b b2a b1b b1a
+ b2b b2a b1a b1b b1a b3b b3a b1b b1a b2a b2b b1a vdd b1b b5b vss vss b2b b1a vdd
+ b0a b0b b0a vdd b0b b0a b0b vss b1a b0a b4a vdd b0b vdd vss b0a b0b vss b1b b0a
+ dac_3v_column_0/dum0_in b0b b0b b0a vdd b0a b0b vdd b0a b0b vdd b2b b3a vdd b0b
+ b0a b0b b0a vdd vdd b0b vss vdd vdd b0a b1a vdd vdd vss vdd b0b m1_6304_841# vdd
+ b0a b0b b3b m1_6304_841# b5a b0a b1b b0b dac_3v_column_dummy
Xdac_3v_column_dummy_1 m1_25325_837# b0a vdd b0b b1b b0a vdd b2a vss vss b4b b1b b2a
+ b1b b1a b2b b2a b1a b1b b1a b3b b3a b1b b1a b2a b2b b1a vdd b1b b5b vss vss b2b
+ b1a vdd b0a b0b b0a vdd b0b b0a b0b vss b1a b0a b4a vdd b0b vdd vss b0a b0b vss
+ b1b b0a m1_25325_837# b0b b0b b0a vdd b0a b0b vdd b0a b0b vdd b2b b3a vdd b0b b0a
+ b0b b0a vdd vdd b0b vss vdd vdd b0a b1a vdd vdd vss vdd b0b Vlow vdd b0a b0b b3b
+ dac_3v_column_odd_7/dum_out1 b5a b0a b1b b0b dac_3v_column_dummy
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0 a_n242_n264# a_50_n42# a_n108_n42#
+ a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n242_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0 a_50_n42# a_n50_n139# w_n308_n339#
+ a_n108_n42#
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n308_n339# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_L7BSKG__0 a_n73_n11# a_n33_n99# a_15_n11# a_n175_n185#
X0 a_15_n11# a_n33_n99# a_n73_n11# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_LGS3BL__0 a_n73_n64# a_n33_n161# a_15_n64# w_n211_n284#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n211_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_64Z3AY__0 a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt rc_osc_level_shifter__0 out_h outb_h in_l inb_l avss dvdd avdd dvss
XXM15 outb_h out_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM16 avdd outb_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM17 avss outb_h avss in_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM18 avss avss out_h inb_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM19 m1_2204_n1198# out_h avdd avdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM7 dvdd in_l inb_l dvdd sky130_fd_pr__pfet_01v8_LGS3BL__0
XXM8 inb_l dvss in_l dvss sky130_fd_pr__nfet_01v8_64Z3AY__0
XXM20 m1_2204_n1198# outb_h avdd out_h sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ a_n2110_1084# a_2206_1084# a_1708_n1516#
+ a_4696_1084# a_48_1084# a_n2442_n1516# a_n1612_1084# a_n4600_1084# a_1708_1084#
+ a_3202_n1516# a_n1446_n1516# a_2870_1084# a_712_1084# a_n284_n1516# a_4696_n1516#
+ a_5028_1084# a_n948_1084# a_2206_n1516# a_n1446_1084# a_n4434_1084# a_n616_n1516#
+ a_3202_1084# a_546_1084# a_1210_n1516# a_n3936_1084# a_5194_n1516# a_2704_1084#
+ a_n4766_n1516# a_n4268_1084# a_3036_1084# a_4198_n1516# a_5526_n1516# a_878_n1516#
+ a_n118_n1516# a_n2442_1084# a_n3770_n1516# a_n5430_1084# a_2538_1084# a_1210_1084#
+ a_5526_1084# a_n5264_n1516# a_4530_n1516# a_n2774_n1516# a_n1944_1084# a_n4932_1084#
+ a_n450_1084# a_n4268_n1516# a_3700_1084# a_3534_n1516# a_n1778_n1516# a_n2276_1084#
+ a_5028_n1516# a_n5264_1084# a_1044_1084# a_4032_1084# a_2538_n1516# a_n3272_n1516#
+ a_n1778_1084# a_n4600_n1516# a_n4766_1084# a_n284_1084# a_n948_n1516# a_3534_1084#
+ a_380_n1516# a_878_1084# a_4032_n1516# a_n2276_n1516# a_n3604_n1516# a_n5098_1084#
+ a_n2940_1084# a_1542_n1516# a_712_n1516# a_3036_n1516# a_n2608_n1516# a_n3272_1084#
+ a_3368_1084# a_2040_1084# a_n1280_n1516# a_n118_1084# a_n4102_n1516# a_n2774_1084#
+ a_2040_n1516# a_1542_1084# a_4530_1084# a_n1612_n1516# a_n5596_n1516# a_4862_n1516#
+ a_n450_n1516# a_n3106_n1516# a_1044_n1516# a_n782_1084# a_214_n1516# a_n3106_1084#
+ a_3866_n1516# a_n5596_1084# a_n1280_1084# a_1376_1084# a_4364_1084# a_n2110_n1516#
+ a_n5726_n1646# a_n2608_1084# a_380_1084# a_5360_n1516# a_n3770_1084# a_n4932_n1516#
+ a_3866_1084# a_n1114_n1516# a_2870_n1516# a_n5098_n1516# a_4364_n1516# a_n616_1084#
+ a_n3936_n1516# a_1874_n1516# a_4198_1084# a_3368_n1516# a_n1114_1084# a_n4102_1084#
+ a_48_n1516# a_n5430_n1516# a_2372_1084# a_5360_1084# a_214_1084# a_n2940_n1516#
+ a_n3604_1084# a_n4434_n1516# a_1874_1084# a_2372_n1516# a_3700_n1516# a_4862_1084#
+ a_n1944_n1516# a_n3438_n1516# a_n782_n1516# a_1376_n1516# a_2704_n1516# a_5194_1084#
+ a_546_n1516# a_n3438_1084#
X0 a_n4932_1084# a_n4932_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X1 a_1376_1084# a_1376_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X2 a_878_1084# a_878_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X3 a_4198_1084# a_4198_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X4 a_3700_1084# a_3700_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X5 a_n3770_1084# a_n3770_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X6 a_n1446_1084# a_n1446_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X7 a_n4268_1084# a_n4268_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X8 a_n2110_1084# a_n2110_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X9 a_1874_1084# a_1874_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X10 a_2372_1084# a_2372_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X11 a_2538_1084# a_2538_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X12 a_4696_1084# a_4696_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X13 a_3036_1084# a_3036_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X14 a_5194_1084# a_5194_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X15 a_n1944_1084# a_n1944_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X16 a_n4766_1084# a_n4766_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X17 a_n2608_1084# a_n2608_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X18 a_n2442_1084# a_n2442_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X19 a_214_1084# a_214_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X20 a_n5430_1084# a_n5430_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X21 a_n5264_1084# a_n5264_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X22 a_n3106_1084# a_n3106_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X23 a_2870_1084# a_2870_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X24 a_n1280_1084# a_n1280_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X25 a_1210_1084# a_1210_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X26 a_3534_1084# a_3534_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X27 a_712_1084# a_712_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X28 a_4032_1084# a_4032_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X29 a_n118_1084# a_n118_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X30 a_n3604_1084# a_n3604_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X31 a_n4102_1084# a_n4102_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X32 a_n1778_1084# a_n1778_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X33 a_n4600_1084# a_n4600_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X34 a_n2276_1084# a_n2276_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X35 a_4530_1084# a_4530_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X36 a_n5098_1084# a_n5098_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X37 a_n616_1084# a_n616_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X38 a_1044_1084# a_1044_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X39 a_3368_1084# a_3368_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X40 a_380_1084# a_380_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X41 a_546_1084# a_546_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X42 a_n2940_1084# a_n2940_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X43 a_n2774_1084# a_n2774_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X44 a_n5596_1084# a_n5596_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X45 a_n3438_1084# a_n3438_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X46 a_n3272_1084# a_n3272_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X47 a_n1114_1084# a_n1114_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X48 a_1542_1084# a_1542_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X49 a_1708_1084# a_1708_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X50 a_3866_1084# a_3866_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X51 a_2040_1084# a_2040_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X52 a_2206_1084# a_2206_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X53 a_4364_1084# a_4364_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X54 a_5028_1084# a_5028_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X55 a_n3936_1084# a_n3936_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X56 a_n450_1084# a_n450_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X57 a_n284_1084# a_n284_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X58 a_n4434_1084# a_n4434_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X59 a_n1612_1084# a_n1612_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X60 a_48_1084# a_48_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X61 a_2704_1084# a_2704_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X62 a_4862_1084# a_4862_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X63 a_3202_1084# a_3202_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X64 a_5360_1084# a_5360_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X65 a_5526_1084# a_5526_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X66 a_n948_1084# a_n948_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
X67 a_n782_1084# a_n782_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=11
.ends

.subckt sky130_fd_pr__nfet_01v8_L9WNCD__0 a_15_n19# a_n175_n193# a_n73_n19# a_n33_n107#
X0 a_15_n19# a_n33_n107# a_n73_n19# a_n175_n193# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__2 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_AZFCP3 m3_n486_n640# c1_n446_n600#
X0 c1_n446_n600# m3_n486_n640# sky130_fd_pr__cap_mim_m3_1 l=6 w=3
.ends

.subckt sky130_fd_pr__pfet_01v8_2Z69BZ__0 w_n211_n226# a_n73_n6# a_15_n6# a_n33_n103#
X0 a_15_n6# a_n33_n103# a_n73_n6# w_n211_n226# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_ef_ip__rc_osc_500k avdd dvdd ena dout dvss avss
XXM12 avss m1_7544_4585# avss m1_2993_5163# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM23 avss m1_6353_4130# m1_513_6590# rc_osc_level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM34 avdd rc_osc_level_shifter_0/out_h avdd m1_2336_4786# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM13 avss m1_7758_4785# m1_7544_4585# ena sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM24 avdd m1_2336_4786# avdd m1_2985_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM25 avdd m1_2336_4786# avdd m1_3601_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM35 dout rc_osc_level_shifter_0/inb_l dvss dvss sky130_fd_pr__nfet_01v8_L7BSKG__0
XXM36 avss m1_2561_4188# m1_2336_4786# rc_osc_level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM15 m1_5347_4782# m1_4789_4781# avdd m1_5449_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM26 avdd m1_2336_4786# avdd m1_4217_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM37 m1_2993_5163# m1_5910_4786# avdd m1_6681_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM16 avss m1_5347_4782# m1_5128_4639# m1_4789_4781# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM27 avss m1_4016_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM38 avss m1_2993_5163# m1_6240_4639# m1_5910_4786# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM17 avdd m1_2336_4786# avdd m1_4833_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM28 avss m1_3460_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM39 avdd m1_2336_4786# avdd m1_6065_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
Xrc_osc_level_shifter_0 rc_osc_level_shifter_0/out_h rc_osc_level_shifter_0/outb_h
+ ena rc_osc_level_shifter_0/inb_l avss dvdd avdd dvss rc_osc_level_shifter__0
XXM18 avdd m1_2336_4786# avdd m1_5449_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM29 avss m1_2904_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM19 avss m1_5128_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
Xsky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_0 avdd m1_8336_3118# m1_7838_518# m1_10660_3118#
+ m1_6012_3118# avdd m1_4352_3118# avdd m1_7672_3118# m1_9166_518# m1_4518_518# m1_9000_3118#
+ m1_6676_3118# m1_5846_518# m1_10826_518# m1_10992_3118# m1_5016_3118# m1_8170_518#
+ m1_4684_3118# avdd m1_5514_518# m1_9332_3118# m1_6676_3118# m1_7174_518# avdd m1_11158_518#
+ m1_8668_3118# avdd avdd m1_9000_3118# m1_10162_518# m1_11490_518# m1_6842_518# m1_5846_518#
+ avdd avdd avdd m1_8668_3118# m1_7340_3118# m1_10494_4056# avdd m1_10494_518# avdd
+ avdd avdd m1_5680_3118# avdd m1_9664_3118# m1_9498_518# m1_4186_518# avdd m1_11158_518#
+ avdd m1_7008_3118# m1_9996_3118# m1_8502_518# avdd m1_4352_3118# avdd avdd m1_5680_3118#
+ m1_5182_518# m1_9664_3118# m1_6510_518# m1_7008_3118# m1_10162_518# avdd avdd avdd
+ avdd m1_7506_518# m1_6842_518# m1_9166_518# avdd avdd m1_9332_3118# m1_8004_3118#
+ m1_4850_518# m1_6012_3118# avdd avdd m1_8170_518# m1_7672_3118# m1_10660_3118# m1_4518_518#
+ avdd m1_10826_518# m1_5514_518# avdd m1_7174_518# m1_5348_3118# m1_6178_518# avdd
+ m1_9830_518# avdd m1_4684_3118# m1_7340_3118# m1_10328_3118# avdd avss avdd m1_6344_3118#
+ m1_11490_518# avdd avdd m1_9996_3118# m1_4850_518# m1_8834_518# avdd m1_10494_518#
+ m1_5348_3118# avdd m1_7838_518# m1_10328_3118# m1_9498_518# m1_5016_3118# avdd m1_6178_518#
+ avdd m1_8336_3118# m1_11324_3118# m1_6344_3118# avdd avdd avdd m1_8004_3118# m1_8502_518#
+ m1_9830_518# m1_10992_3118# m1_4186_518# avdd m1_5182_518# m1_7506_518# m1_8834_518#
+ m1_11324_3118# m1_6510_518# avdd sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ
Xsky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_1 m1_3834_9768# m1_8150_9768# m1_7652_7168#
+ m1_10806_9768# m1_6158_9768# m1_3668_7168# m1_4498_9768# m1_1510_9768# m1_7818_9768#
+ m1_9312_7168# m1_4664_7168# m1_8814_9768# m1_6822_9768# m1_5660_7168# m1_10640_7168#
+ m1_11138_9768# m1_5162_9768# m1_8316_7168# m1_4498_9768# m1_1510_9768# m1_5328_7168#
+ m1_9146_9768# m1_6490_9768# m1_7320_7168# m1_2174_9768# m1_11304_7168# m1_8814_9768#
+ m1_1344_7168# m1_1842_9768# m1_9146_9768# m1_10308_7168# m1_10494_4056# m1_6988_7168#
+ m1_5992_7168# m1_3502_9768# m1_2340_7168# m1_514_9768# m1_8482_9768# m1_7154_9768#
+ m1_11470_9768# m1_680_7168# m1_10640_7168# m1_3336_7168# m1_4166_9768# m1_1178_9768#
+ m1_5494_9768# m1_1676_7168# m1_9810_9768# m1_9644_7168# m1_4332_7168# m1_3834_9768#
+ m1_10972_7168# m1_846_9768# m1_7154_9768# m1_10142_9768# m1_8648_7168# m1_2672_7168#
+ m1_4166_9768# m1_1344_7168# m1_1178_9768# m1_5826_9768# m1_4996_7168# m1_9478_9768#
+ m1_6324_7168# m1_6822_9768# m1_9976_7168# m1_3668_7168# m1_2340_7168# m1_846_9768#
+ m1_3170_9768# m1_7652_7168# m1_6656_7168# m1_8980_7168# m1_3336_7168# m1_2838_9768#
+ m1_9478_9768# m1_8150_9768# m1_4664_7168# m1_5826_9768# m1_2008_7168# m1_3170_9768#
+ m1_7984_7168# m1_7486_9768# m1_10474_9768# m1_4332_7168# m1_513_6590# m1_10972_7168#
+ m1_5660_7168# m1_3004_7168# m1_6988_7168# m1_5162_9768# m1_6324_7168# m1_2838_9768#
+ m1_9976_7168# m1_514_9768# m1_4830_9768# m1_7486_9768# m1_10474_9768# m1_4000_7168#
+ avss m1_3502_9768# m1_6490_9768# m1_11304_7168# m1_2174_9768# m1_1012_7168# m1_9810_9768#
+ m1_4996_7168# m1_8980_7168# m1_1012_7168# m1_10308_7168# m1_5494_9768# m1_2008_7168#
+ m1_7984_7168# m1_10142_9768# m1_9312_7168# m1_4830_9768# m1_1842_9768# m1_5992_7168#
+ m1_680_7168# m1_8482_9768# m1_11470_9768# m1_6158_9768# m1_3004_7168# m1_2506_9768#
+ m1_1676_7168# m1_7818_9768# m1_8316_7168# m1_9644_7168# m1_10806_9768# m1_4000_7168#
+ m1_2672_7168# m1_5328_7168# m1_7320_7168# m1_8648_7168# m1_11138_9768# m1_6656_7168#
+ m1_2506_9768# sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ
XXM1 avss m1_3128_4787# m1_2904_4639# m1_2993_5163# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM2 m1_3128_4787# m1_2993_5163# avdd m1_2985_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM3 m1_3679_4781# m1_3128_4787# avdd m1_3601_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM4 avss m1_3679_4781# m1_3460_4639# m1_3128_4787# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
Xsky130_fd_pr__nfet_01v8_L9WNCD_0 m1_11938_5890# dvss dvss m1_7758_4785# sky130_fd_pr__nfet_01v8_L9WNCD__0
XXM5 m1_11938_5890# dvss dout ena sky130_fd_pr__nfet_01v8_L9WNCD__0
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__2
XXM7 m1_4789_4781# m1_4235_4789# avdd m1_4833_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM8 avss m1_4789_4781# m1_4572_4639# m1_4235_4789# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM9 m1_4235_4789# m1_3679_4781# avdd m1_4217_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
Xsky130_fd_pr__pfet_01v8_LGS3BL_0 dvdd m1_7758_4785# dout dvdd sky130_fd_pr__pfet_01v8_LGS3BL__0
XXC1 avss m1_3128_4787# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC2 avss m1_3679_4781# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC3 avss m1_4235_4789# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC4 avss m1_4789_4781# sky130_fd_pr__cap_mim_m3_1_AZFCP3
Xsky130_fd_pr__pfet_01v8_2Z69BZ_0 dvdd m1_7758_4785# dvdd ena sky130_fd_pr__pfet_01v8_2Z69BZ__0
Xsky130_fd_pr__cap_mim_m3_1_AZFCP3_1 avss m1_5347_4782# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXM40 avdd m1_2336_4786# avdd m1_6681_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM30 avss m1_2561_4188# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM41 avss m1_6240_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM20 avss m1_4572_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM31 m1_5910_4786# m1_5347_4782# avdd m1_6065_5653# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM42 avss m1_5684_4639# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM10 avss m1_4235_4789# m1_4016_4639# m1_3679_4781# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM21 avss m1_6353_4130# avss m1_6353_4130# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM32 avss m1_5910_4786# m1_5684_4639# m1_5347_4782# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
XXM11 m1_7758_4785# m1_2993_5163# avdd dvdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM22 avdd m1_2336_4786# avdd m1_2336_4786# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH__0
XXM33 avss m1_6353_4130# avss rc_osc_level_shifter_0/outb_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR__0
.ends

.subckt chipalooza_testchip_2 gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17]
+ gpio_analog[1] gpio_analog[5] gpio_analog[6] gpio_analog[8] gpio_analog[9] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[7] io_analog[0] io_analog[10] io_analog[1]
+ io_analog[2] io_analog[3] io_analog[4] io_analog[7] io_analog[8] io_analog[9] io_analog[5]
+ io_analog[6] io_oeb[0] io_oeb[12] io_oeb[13] io_oeb[17] io_oeb[1] io_oeb[23] io_oeb[24]
+ io_oeb[25] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_out[0] io_out[12] io_out[13] io_out[17] io_out[1] io_out[23] io_out[24] io_out[25]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[120] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[11] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65]
+ la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70]
+ la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75]
+ la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80]
+ la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85]
+ la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90]
+ la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95]
+ la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] vccd1
+ vccd2 vdda1 vdda2 sky130_aa_ip__programmable_pll_0/D10 sky130_aa_ip__programmable_pll_0/S4
+ m2_35602_800# power_stage_1[2]/p_in ct2_switch_array_1/switch_array_2_0/channel0_in_to_out[0]
+ m3_800_35586# m3_800_463198# sky130_aa_ip__programmable_pll_0/S1 sky130_aa_ip__programmable_pll_0/D13
+ sky130_ef_ip__idac3v_8bit_0/din[0] m2_106522_800# sky130_ef_ip__rheostat_8bit_0/b1
+ power_stage_0[1]/p_in ct2_switch_array_10/switch_array_2_0/channel0_in_to_out[1]
+ ct2_switch_array_9/switch_array_2_0/channel1_out m2_335830_800# m2_86428_800# m3_584320_272394#
+ m2_58060_800# m3_800_512330# power_stage_1[6]/p_in ct2_switch_array_4/switch_array_2_0/channel0_in_to_out[0]
+ m3_800_508784# ct2_switch_array_4/switch_array_2_0/channel1_out m2_29692_800# m2_40330_800#
+ m2_11962_800# ct2_switch_array_12/switch_array_2_0/channel1_out sky130_ef_ip__rheostat_8bit_0/b4
+ m2_403204_800# sky130_aa_ip__programmable_pll_0/D5 m2_111250_800# m2_28510_800#
+ sky130_ef_ip__rdac3v_8bit_0/b7 m3_800_466744# m3_800_506420# power_stage_0[6]/p_in
+ sky130_ef_ip__cdac3v_12bit_0/SELD0 m3_584320_7072# sky130_ef_ip__idac3v_8bit_0/din[3]
+ m2_91156_800# sky130_aa_ip__programmable_pll_0/S5 sky130_ef_ip__rheostat_8bit_0/b6
+ m3_584318_93554# m2_62788_800# m2_268456_800# m4_319794_703100# ct2_switch_array_3/switch_array_2_0/channel0_in_to_out[1]
+ m3_584288_359674# m2_79336_800# m2_430390_800# m3_584000_412006# m2_7234_800# sky130_ef_ip__idac3v_8bit_0/din[7]
+ m2_391384_800# m2_61606_800# m3_584180_92372# m4_176694_703100# ct2_switch_array_11/switch_array_2_0/channel0_in_to_out[1]
+ ct2_switch_array_8/switch_array_2_0/channel1_in_to_out[0] m3_800_249652# m3_800_5890#
+ ct2_switch_array_13/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_5/switch_array_2_0/channel1_in_to_out[1]
+ m2_357106_800# sky130_aa_ip__programmable_pll_0/DN_INPUT ct2_switch_array_9/switch_array_2_0/channel0_in_to_out[1]
+ ct2_switch_array_13/switch_array_2_0/channel1_in_to_out[0] m2_84064_800# ct2_switch_array_6/switch_array_2_0/channel1_in_to_out[0]
+ m2_328738_800# m2_55696_800# power_stage_0[0]/p_in m3_584320_587908# sky130_aa_ip__programmable_pll_0/D17
+ m2_33238_800# power_stage_0[2]/p_in sky130_aa_ip__programmable_pll_0/D9 m2_76972_800#
+ m2_384292_800# m2_4870_800# m2_54514_800# sky130_ef_ip__idac3v_8bit_0/din[1] m3_327594_703100#
+ m2_104158_800# m2_264910_800# ct2_switch_array_2/switch_array_2_0/channel0_in_to_out[1]
+ m3_584320_452882# ct2_switch_array_8/switch_array_2_0/channel1_out m2_125434_800#
+ sky130_aa_ip__programmable_pll_0/OUT sky130_aa_ip__programmable_pll_0/S7 ct2_switch_array_0/switch_array_2_0/channel0_in_to_out[0]
+ ct2_switch_array_13/switch_array_2_0/channel0_in_to_out[0] sky130_ef_ip__idac3v_8bit_0/ref_sel_vbg
+ ct2_switch_array_10/switch_array_2_0/channel1_in_to_out[1] m3_584320_12982# m2_423298_800#
+ sky130_ef_ip__rheostat_8bit_0/b5 m3_800_122030# power_stage_1[4]/p_in m2_26146_800#
+ m2_444574_800# sky130_ef_ip__samplehold_0/ena m2_30874_800# m2_69880_800# m3_800_335896#
+ sky130_ef_ip__cdac3v_12bit_0/SELD11 m2_47422_800# ct2_switch_array_4/switch_array_2_0/channel1_in_to_out[0]
+ m3_584320_406096# m2_101794_800# m4_228394_703100# m3_800_77626# ct2_switch_array_3/switch_array_2_0/channel1_out
+ m2_584050_800# sky130_ak_ip__cmos_vref_0/trim3 m2_118342_800# ct2_switch_array_7/switch_array_2_0/channel1_out
+ m3_800_293856# ct2_switch_array_8/switch_array_2_0/channel0_in_to_out[0] sky130_ak_ip__cmos_vref_0/trim2
+ m3_800_333532# sky130_ef_ip__rdac3v_8bit_0/b0 ct2_switch_array_15/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__cdac3v_12bit_0/SELD9 m2_100612_800# m2_98248_800# m2_80518_800# m2_52150_800#
+ ct2_switch_array_15/switch_array_2_0/channel1_in_to_out[1] sky130_aa_ip__programmable_pll_0/S6
+ ct2_switch_array_3/switch_array_2_0/channel1_in_to_out[1] m2_19054_800# m3_584318_48896#
+ m2_437482_800# m2_257818_800# m2_23782_800# ct2_switch_array_7/switch_array_2_0/channel0_in_to_out[0]
+ m3_800_2344# m3_584320_409642# sky130_aa_ip__programmable_pll_0/D15 m2_398476_800#
+ m3_800_14164# m2_123070_800# m2_292096_800# ct2_switch_array_9/switch_array_2_0/channel1_in_to_out[0]
+ m2_380746_800# ct2_switch_array_10/switch_array_2_0/channel1_out m2_22600_800# sky130_aa_ip__programmable_pll_0/OUTB
+ sky130_am_ip__ldo_01v8_0/ENA ct2_switch_array_12/switch_array_2_0/channel0_in_to_out[0]
+ m3_584316_22438# m2_95884_800# power_stage_0[5]/p_in m2_73426_800# m2_1324_800#
+ m5_319794_703100# m3_584320_497304# ct2_switch_array_6/switch_array_2_0/channel0_in_to_out[1]
+ m2_16690_800# m2_94702_800# m4_166394_703100# m2_352378_800# m2_412660_800# m2_581686_800#
+ m2_373654_800# m2_115978_800# m5_176694_703100# sky130_aa_ip__programmable_pll_0/PRE_SCALAR
+ ct2_switch_array_2/switch_array_2_0/channel1_in_to_out[1] m2_394930_800# m3_171694_703100#
+ ct2_switch_array_0/switch_array_2_0/channel1_out m2_580504_800# ct2_switch_array_0/switch_array_2_0/channel1_in_to_out[0]
+ m2_45058_800# ct2_switch_array_14/switch_array_2_0/channel1_in_to_out[1] m3_584112_456428#
+ m2_88792_800# m2_441028_800# m2_66334_800# sky130_aa_ip__programmable_pll_0/OUT_CORE
+ m2_37966_800# sky130_ef_ip__rdac3v_8bit_0/b6 m2_87610_800# sky130_ef_ip__rdac3v_8bit_0/b4
+ m2_345286_800# sky130_ef_ip__cdac3v_12bit_0/SELD1 m2_15508_800# m2_433936_800# sky130_ef_ip__cdac3v_12bit_0/SELD6
+ m2_574594_800# m2_366562_800# m2_108886_800# sky130_aa_ip__programmable_pll_0/D0
+ m3_800_423522# m3_584320_316816# m2_260182_800# m3_174194_703100# m3_800_419976#
+ m3_584320_365584# m2_71062_800# m2_107704_800# ct2_switch_array_1/switch_array_2_0/channel0_in_to_out[1]
+ sky130_icrg_ip__ulpcomp2_0/vout ct2_switch_array_1/switch_array_2_0/channel1_out
+ m2_42694_800# m3_800_465562# m2_20236_800# m2_59242_800# sky130_aa_ip__programmable_pll_0/DIV_OUT
+ m2_63970_800# m2_405568_800# m3_584320_363220# ct2_switch_array_11/switch_array_2_0/channel1_in_to_out[0]
+ m3_584320_454064# m2_371290_800# m2_41512_800# m3_800_16528# m3_800_79990# m2_338194_800#
+ sky130_aa_ip__programmable_pll_0/S2 ct2_switch_array_7/switch_array_2_0/channel1_in_to_out[0]
+ m4_218094_703100# m2_426844_800# m2_299188_800# m2_320464_800# m2_387838_800# m2_359470_800#
+ m2_112432_800# m2_281458_800# m5_228394_703100# ct2_switch_array_5/switch_array_2_0/channel0_in_to_out[0]
+ m2_341740_800# m2_92338_800# ct2_switch_array_12/switch_array_2_0/channel1_in_to_out[0]
+ m2_9598_800# sky130_aa_ip__programmable_pll_0/D14 sky130_ef_ip__idac3v_8bit_0/din[5]
+ m2_410296_800# m3_223394_703100# ct2_switch_array_13/switch_array_2_0/channel1_in_to_out[1]
+ m3_800_337078# ct2_switch_array_10/switch_array_2_0/channel1_in_to_out[0] sky130_ef_ip__rheostat_8bit_0/b3
+ m3_584320_3526# sky130_ef_ip__idac3v_8bit_0/ena m2_13144_800# m2_431572_800# m2_8416_800#
+ ct2_switch_array_1/switch_array_2_0/channel1_in_to_out[1] ct2_switch_array_11/switch_array_2_0/channel1_out
+ m2_392566_800# ct2_switch_array_12/switch_array_2_0/channel0_in_to_out[1] sky130_ef_ip__rc_osc_500k_1/ena
+ m2_34420_800# sky130_aa_ip__programmable_pll_0/D8 ct2_switch_array_2/switch_array_2_0/channel1_out
+ m2_370108_800# ct2_switch_array_6/switch_array_2_0/channel1_in_to_out[1] sky130_ef_ip__rdac3v_8bit_0/b1
+ m3_584320_586726# m2_419752_800# sky130_ef_ip__samplehold_0/hold sky130_ef_ip__cdac3v_12bit_0/SELD10
+ m2_313372_800# m2_105340_800# sky130_aa_ip__programmable_pll_0/D12 sky130_ak_ip__cmos_vref_0/trim1
+ m2_274366_800# li_477734_350840# m2_542680_800# m2_85246_800# sky130_ef_ip__cdac3v_12bit_0/RST
+ sky130_ef_ip__rc_osc_16M_0/dout m2_295642_800# m2_56878_800# m2_364198_800# ct2_switch_array_9/switch_array_2_0/channel0_in_to_out[0]
+ m3_800_36768# m2_424480_800# sky130_ef_ip__idac3v_8bit_0/din[6] m2_10780_800# ct2_switch_array_0/switch_array_2_0/channel0_in_to_out[1]
+ m4_330094_703100# sky130_aa_ip__programmable_pll_0/D3 sky130_ef_ip__rheostat_8bit_0/b2
+ sky130_iic_ip__audiodac_drv_lite_0/in_p m2_385474_800# m2_402022_800# power_stage_0[4]/p_in
+ m2_127798_800# m2_363016_800# m3_584320_362038# ct2_switch_array_8/switch_array_2_0/channel1_in_to_out[1]
+ m3_584320_273576# m5_166394_703100# power_stage_1[1]/p_in m2_334648_800# m3_800_509966#
+ m2_306280_800# m2_267274_800# sky130_aa_ip__programmable_pll_0/D1 m2_355924_800#
+ ct2_switch_array_14/switch_array_2_0/channel1_out m2_78154_800# m2_82882_800# m2_288550_800#
+ ct2_switch_array_4/switch_array_2_0/channel1_in_to_out[1] m2_6052_800# sky130_icrg_ip__ulpcomp2_0/clk
+ m3_800_76444# ct2_switch_array_5/switch_array_2_0/channel1_out m2_49786_800# m2_60424_800#
+ m2_99430_800# sky130_am_ip__ldo_01v8_0/SEL_EXT m3_800_292674# sky130_ef_ip__idac3v_8bit_0/din[2]
+ m2_110068_800# m2_270820_800# m3_584320_8254# m2_27328_800# m3_800_247288# ct2_switch_array_3/switch_array_2_0/channel0_in_to_out[0]
+ m2_445756_800# sky130_ef_ip__ccomp3v_cl_0/ENA sky130_ef_ip__rheostat_8bit_0/b7 ct2_switch_array_8/switch_array_2_0/channel0_in_to_out[1]
+ m2_81700_800# m2_378382_800# m2_48604_800# m3_583898_21256# m2_360652_800# m2_102976_800#
+ m3_800_290310# sky130_ef_ip__cdac3v_12bit_0/SELD3 m2_327556_800# m3_584320_408460#
+ m2_377200_800# sky130_ef_ip__rheostat_8bit_0/b0 m2_119524_800# sky130_aa_ip__programmable_pll_0/S3
+ ct2_switch_array_11/switch_array_2_0/channel1_in_to_out[1] ct2_switch_array_7/switch_array_2_0/channel0_in_to_out[1]
+ m2_348832_800# m2_32056_800# ct2_switch_array_5/switch_array_2_0/channel1_in_to_out[0]
+ sky130_aa_ip__programmable_pll_0/OUT_USB m2_75790_800# m2_417388_800# m2_53332_800#
+ sky130_ef_ip__cdac3v_12bit_0/SELD2 sky130_ef_ip__rdac3v_8bit_0/ena m3_584320_498486#
+ m3_584288_364404# sky130_aa_ip__programmable_pll_0/UP_INPUT m2_438664_800# sky130_aa_ip__programmable_pll_0/D19
+ m2_24964_800# m2_332284_800# m2_399658_800# m2_416206_800# m2_124252_800# sky130_aa_ip__programmable_pll_0/UP_OUT
+ m2_420934_800# m2_212902_800# ct2_switch_array_4/switch_array_2_0/channel0_in_to_out[1]
+ power_stage_1[0]/p_in sky130_ak_ip__cmos_vref_0/trim0 m2_381928_800# m2_353560_800#
+ m2_578140_800# m5_218094_703100# m2_331102_800# m3_800_10618# sky130_ef_ip__cdac3v_12bit_0/SELD7
+ ct2_switch_array_2/switch_array_2_0/channel0_in_to_out[0] sky130_aa_ip__programmable_pll_0/D4
+ m3_800_379118# m2_549772_800# m2_3688_800# m2_302734_800# sky130_ef_ip__rdac3v_8bit_0/b2
+ sky130_ef_ip__cdac3v_12bit_0/SELD4 m3_325094_703100# m2_263728_800# m2_74608_800#
+ m2_46240_800# m2_2506_800# sky130_ef_ip__cdac3v_12bit_0/SELD5 sky130_ef_ip__rdac3v_8bit_0/b5
+ m2_442210_800# m2_17872_800# m2_325192_800# m2_409114_800# m2_117160_800# ct2_switch_array_0/switch_array_2_0/channel1_in_to_out[1]
+ m3_800_123212# ct2_switch_array_3/switch_array_2_0/channel1_in_to_out[0] m2_413842_800#
+ m2_582868_800# sky130_ef_ip__idac3v_8bit_0/din[4] m3_800_119666# m2_374836_800#
+ sky130_iic_ip__audiodac_drv_lite_0/in_n m3_319794_703100# power_stage_1[3]/p_in
+ m3_584320_317998# m2_97066_800# sky130_icrg_ip__ulpcomp2_0/ena sky130_ak_ip__cmos_vref_0/ena
+ m2_324010_800# m2_68698_800# m3_584320_11800# m2_285004_800# m3_583600_16528# sky130_aa_ip__programmable_pll_0/D18
+ m3_176694_703100# m3_800_78808# m2_50968_800# m2_256636_800# m2_89974_800# ct2_switch_array_9/switch_array_2_0/channel1_in_to_out[1]
+ m3_800_422340# m2_67516_800# sky130_aa_ip__programmable_pll_0/D16 m2_277912_800#
+ sky130_ef_ip__rdac3v_8bit_0/b3 m2_121888_800# ct2_switch_array_1/switch_array_2_0/channel1_in_to_out[0]
+ m2_346468_800# m2_396112_800# m3_800_380300# m5_330094_703100# m3_584318_17710#
+ m2_406750_800# power_stage_1[5]/p_in m2_367744_800# m2_120706_800# sky130_aa_ip__programmable_pll_0/D6
+ power_stage_0[3]/p_in m3_800_3526# m2_553318_800# m2_261364_800# m3_800_15346# ct2_switch_array_11/switch_array_2_0/channel0_in_to_out[0]
+ m2_72244_800# m2_316918_800# sky130_ef_ip__cdac3v_12bit_0/SELD8 m2_39148_800# ct2_switch_array_15/switch_array_2_0/channel0_in_to_out[1]
+ ct2_switch_array_7/switch_array_2_0/channel1_in_to_out[1] m2_43876_800# m2_93520_800#
+ m2_435118_800# m2_21418_800# m3_225894_703100# m3_583894_47714# ct2_switch_array_5/switch_array_2_0/channel0_in_to_out[1]
+ m2_114796_800# m2_339376_800# w_533663_487548# m2_350014_800# m2_389020_800# ct2_switch_array_6/switch_array_2_0/channel0_in_to_out[0]
+ m3_584320_2344# ct2_switch_array_12/switch_array_2_0/channel1_in_to_out[1] m2_321646_800#
+ m3_584320_450518# m2_113614_800# sky130_ef_ip__rc_osc_16M_0/ena m2_546226_800# sky130_aa_ip__programmable_pll_0/D7
+ m2_254272_800# m3_800_250834# ct2_switch_array_14/switch_array_2_0/channel0_in_to_out[1]
+ m2_342922_800# m2_65152_800# m2_309826_800# ct2_switch_array_2/switch_array_2_0/channel1_in_to_out[0]
+ vssd1 vssd2 m2_36784_800# sky130_aa_ip__programmable_pll_0/D2 m3_1168_469108# vssa2
+ vssa1 m2_428026_800# m3_228394_703100# m2_14326_800#
Xsky130_ef_ip__rc_osc_16M_0 io_analog[6] vccd2 sky130_ef_ip__rc_osc_16M_0/ena sky130_ef_ip__rc_osc_16M_0/dout
+ vssd2 vssa2 sky130_ef_ip__rc_osc_16M
Xpower_stage_0[0] power_stage_0[0]/p_in io_analog[5] vccd2 vccd2 vssd2 vssd2 power_stage
Xpower_stage_0[1] power_stage_0[1]/p_in io_analog[6] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[2] power_stage_0[2]/p_in io_analog[7] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[3] power_stage_0[3]/p_in io_analog[8] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[4] power_stage_0[4]/p_in io_analog[9] vccd2 vccd2 vssd2 vssd2 power_stage
Xpower_stage_0[5] power_stage_0[5]/p_in io_analog[10] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[6] power_stage_0[6]/p_in power_stage_0[6]/sw_node vdda2 vccd2 vssa2
+ vssd2 power_stage
Xsky130_ef_ip__idac3v_8bit_0 sky130_ef_ip__idac3v_8bit_0/din[6] sky130_ef_ip__idac3v_8bit_0/din[3]
+ sky130_ef_ip__idac3v_8bit_0/din[2] sky130_ef_ip__idac3v_8bit_0/din[0] sky130_ef_ip__idac3v_8bit_0/din[1]
+ sky130_ef_ip__idac3v_8bit_0/din[5] sky130_ef_ip__idac3v_8bit_0/din[4] sky130_ef_ip__idac3v_8bit_0/din[7]
+ sky130_ef_ip__idac3v_8bit_0/ref_sel_vbg sky130_ef_ip__idac3v_8bit_0/ena bias_reference_voltage
+ sky130_ef_ip__idac3v_8bit_0/snk_out sky130_ef_ip__idac3v_8bit_0/src_out sky130_ef_ip__idac3v_8bit_0/ref_in
+ power_stage_0[6]/sw_node vccd2 vssa2 vssd2 sky130_ef_ip__idac3v_8bit
Xpower_stage_1[0] power_stage_1[0]/p_in io_analog[0] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[1] power_stage_1[1]/p_in io_analog[1] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[2] power_stage_1[2]/p_in io_analog[2] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[3] power_stage_1[3]/p_in power_stage_1[3]/sw_node vccd1 vccd1 vssd1
+ vssd1 power_stage
Xpower_stage_1[4] power_stage_1[4]/p_in io_analog[3] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[5] power_stage_1[5]/p_in power_stage_1[5]/sw_node vdda1 vccd1 vssa1
+ vssd1 power_stage
Xpower_stage_1[6] power_stage_1[6]/p_in io_analog[4] vdda1 vccd1 vssa1 vssd1 power_stage
Xsky130_am_ip__ldo_01v8_0 io_analog[10] sky130_am_ip__ldo_01v8_0/VOUT vssa2 sky130_am_ip__ldo_01v8_0/ENA
+ bias_reference_voltage sky130_am_ip__ldo_01v8_0/SEL_EXT vccd2 vssd2 sky130_am_ip__ldo_01v8
Xsky130_ak_ip__cmos_vref_0 sky130_ak_ip__cmos_vref_0/vbg io_analog[9] sky130_ak_ip__cmos_vref_0/ena
+ sky130_ak_ip__cmos_vref_0/vbgsc sky130_ak_ip__cmos_vref_0/vbgtg sky130_ak_ip__cmos_vref_0/trim3
+ sky130_ak_ip__cmos_vref_0/trim2 sky130_ak_ip__cmos_vref_0/trim1 sky130_ak_ip__cmos_vref_0/trim0
+ sky130_ak_ip__cmos_vref_0/vptat vccd2 vssd2 vssd2 sky130_ak_ip__cmos_vref
Xct2_switch_array_0 vccd2 sky130_ef_ip__ccomp3v_cl_0/VINP ct2_switch_array_0/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_0/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_0/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_0/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_0/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__cdac3v_12bit_0/VH vssd2 ct2_switch_array
Xsky130_iic_ip__audiodac_drv_lite_0 sky130_iic_ip__audiodac_drv_lite_0/in_p sky130_iic_ip__audiodac_drv_lite_0/in_n
+ sky130_iic_ip__audiodac_drv_lite_0/out_p sky130_iic_ip__audiodac_drv_lite_0/out_n
+ vccd2 io_analog[5] vssd2 sky130_iic_ip__audiodac_drv_lite
Xsky130_ef_ip__ccomp3v_cl_0 sky130_ef_ip__ccomp3v_cl_0/VINM sky130_ef_ip__ccomp3v_cl_0/VINP
+ io_analog[8] vssa2 vccd2 io_out[17] vssa2 sky130_ef_ip__ccomp3v_cl_0/ENA vssd2 sky130_ef_ip__ccomp3v_cl
Xct2_switch_array_1 vccd2 ct2_switch_array_1/switch_array_2_0/channel0_in ct2_switch_array_1/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_1/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_1/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_1/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_1/switch_array_2_0/channel0_in_to_out[0]
+ sky130_iic_ip__audiodac_drv_lite_0/out_p vssd2 ct2_switch_array
Xsky130_aa_ip__programmable_pll_0 sky130_aa_ip__programmable_pll_0/S6 sky130_aa_ip__programmable_pll_0/UP_INPUT
+ sky130_aa_ip__programmable_pll_0/DN_INPUT sky130_aa_ip__programmable_pll_0/S2 sky130_aa_ip__programmable_pll_0/S3
+ sky130_aa_ip__programmable_pll_0/UP_OUT io_out[12] sky130_aa_ip__programmable_pll_0/ITAIL
+ sky130_aa_ip__programmable_pll_0/S4 sky130_aa_ip__programmable_pll_0/VCTRL_IN sky130_aa_ip__programmable_pll_0/LF_OFFCHIP
+ sky130_aa_ip__programmable_pll_0/S5 sky130_aa_ip__programmable_pll_0/OUT_CORE sky130_aa_ip__programmable_pll_0/OUT_USB
+ sky130_aa_ip__programmable_pll_0/D12 sky130_aa_ip__programmable_pll_0/D13 sky130_aa_ip__programmable_pll_0/D14
+ sky130_aa_ip__programmable_pll_0/D15 sky130_aa_ip__programmable_pll_0/F_IN sky130_aa_ip__programmable_pll_0/D0
+ sky130_aa_ip__programmable_pll_0/D1 sky130_aa_ip__programmable_pll_0/D2 sky130_aa_ip__programmable_pll_0/D3
+ sky130_aa_ip__programmable_pll_0/D4 sky130_aa_ip__programmable_pll_0/D5 sky130_aa_ip__programmable_pll_0/D6
+ sky130_aa_ip__programmable_pll_0/D7 sky130_aa_ip__programmable_pll_0/D8 sky130_aa_ip__programmable_pll_0/D9
+ sky130_aa_ip__programmable_pll_0/D10 sky130_aa_ip__programmable_pll_0/D16 sky130_aa_ip__programmable_pll_0/D17
+ sky130_aa_ip__programmable_pll_0/D18 sky130_aa_ip__programmable_pll_0/D19 sky130_aa_ip__programmable_pll_0/OUTB
+ sky130_aa_ip__programmable_pll_0/OUT sky130_aa_ip__programmable_pll_0/PRE_SCALAR
+ sky130_aa_ip__programmable_pll_0/S1 sky130_aa_ip__programmable_pll_0/S7 sky130_aa_ip__programmable_pll_0/DIV_OUT
+ power_stage_1[3]/sw_node vssd1 sky130_aa_ip__programmable_pll
Xct2_switch_array_2 vccd2 sky130_ef_ip__ccomp3v_cl_0/VINM ct2_switch_array_2/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_2/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_2/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_2/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_2/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__cdac3v_12bit_0/VL vssd2 ct2_switch_array
Xsky130_sw_ip__bgrref_por_0 bias_reference_voltage io_out[7] io_analog[2] vccd1 io_out[8]
+ sky130_sw_ip__bgrref_por_0/porb_h[0] sky130_sw_ip__bgrref_por_0/porb_h[1] vssa1
+ vssd1 sky130_sw_ip__bgrref_por
Xct2_switch_array_3 vccd2 sky130_ef_ip__idac3v_8bit_0/ref_in ct2_switch_array_3/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_3/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_3/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_3/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_3/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ak_ip__cmos_vref_0/vbgtg vssd2 ct2_switch_array
Xct2_switch_array_4 vccd2 sky130_am_ip__ldo_01v8_0/VOUT ct2_switch_array_4/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_4/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_4/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_4/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_4/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ak_ip__cmos_vref_0/vbgsc vssd2 ct2_switch_array
Xsky130_ef_ip__rheostat_8bit_0 sky130_ef_ip__rheostat_8bit_0/b0 sky130_ef_ip__rheostat_8bit_0/b1
+ sky130_ef_ip__rheostat_8bit_0/b2 sky130_ef_ip__rheostat_8bit_0/b3 sky130_ef_ip__rheostat_8bit_0/b4
+ sky130_ef_ip__rheostat_8bit_0/b5 sky130_ef_ip__rheostat_8bit_0/b6 sky130_ef_ip__rheostat_8bit_0/b7
+ sky130_ef_ip__rheostat_8bit_0/out io_analog[1] vccd1 sky130_ef_ip__rheostat_8bit_0/Vhigh
+ sky130_ef_ip__rheostat_8bit_0/Vlow vssa1 vssd1 sky130_ef_ip__rheostat_8bit
Xct2_switch_array_5 vccd2 sky130_ef_ip__idac3v_8bit_0/snk_out ct2_switch_array_5/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_5/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_5/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_5/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_5/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ak_ip__cmos_vref_0/vbg vssd2 ct2_switch_array
Xct2_switch_array_6 vccd2 sky130_ef_ip__idac3v_8bit_0/src_out ct2_switch_array_6/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_6/switch_array_2_0/channel1_in_to_out[0] gpio_noesd[7] vdda2 vssa2
+ ct2_switch_array_6/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_6/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ak_ip__cmos_vref_0/vptat vssd2 ct2_switch_array
Xsky130_ef_ip__samplehold_0 sky130_ef_ip__samplehold_0/out power_stage_1[5]/sw_node
+ sky130_ef_ip__samplehold_0/hold sky130_ef_ip__samplehold_0/in vccd1 sky130_ef_ip__samplehold_0/ena
+ vssa1 vssd1 sky130_ef_ip__samplehold
Xct2_switch_array_7 vccd2 sky130_aa_ip__programmable_pll_0/F_IN ct2_switch_array_7/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_7/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_7/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_7/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_7/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__cdac3v_12bit_0/OUT vssd2 ct2_switch_array
Xct2_switch_array_8 vccd2 sky130_aa_ip__programmable_pll_0/ITAIL ct2_switch_array_8/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_8/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_8/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_8/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_8/switch_array_2_0/channel0_in_to_out[0]
+ ct2_switch_array_8/switch_array_2_0/channel1_in vssd2 ct2_switch_array
Xct2_switch_array_9 vccd2 sky130_aa_ip__programmable_pll_0/VCTRL_IN ct2_switch_array_9/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_9/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_9/switch_array_2_0/channel1_out
+ vdda2 vssa2 ct2_switch_array_9/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_9/switch_array_2_0/channel0_in_to_out[0]
+ sky130_iic_ip__audiodac_drv_lite_0/out_n vssd2 ct2_switch_array
Xct2_switch_array_10 vccd1 sky130_ef_ip__samplehold_0/out ct2_switch_array_10/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_10/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_10/switch_array_2_0/channel1_out
+ vdda1 vssa1 ct2_switch_array_10/switch_array_2_0/channel0_in_to_out[1] la_data_in[117]
+ sky130_icrg_ip__ulpcomp2_0/vinn vssd1 ct2_switch_array
Xct2_switch_array_11 vccd1 sky130_ef_ip__rheostat_8bit_0/out ct2_switch_array_11/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_11/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_11/switch_array_2_0/channel1_out
+ vdda1 vssa1 ct2_switch_array_11/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_11/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__rdac3v_8bit_0/out vssd1 ct2_switch_array
Xsky130_icrg_ip__ulpcomp2_0 sky130_icrg_ip__ulpcomp2_0/ena sky130_icrg_ip__ulpcomp2_0/vout
+ sky130_icrg_ip__ulpcomp2_0/vinn sky130_icrg_ip__ulpcomp2_0/vinp sky130_icrg_ip__ulpcomp2_0/clk
+ vccd1 io_analog[3] vssa1 w_533663_487548# vssd1 sky130_icrg_ip__ulpcomp2
Xct2_switch_array_12 vccd1 sky130_ef_ip__rdac3v_8bit_0/Vlow ct2_switch_array_12/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_12/switch_array_2_0/channel1_in_to_out[0] ct2_switch_array_12/switch_array_2_0/channel1_out
+ vdda1 vssa1 ct2_switch_array_12/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_12/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__rheostat_8bit_0/Vlow vssd1 ct2_switch_array
Xct2_switch_array_13 vccd1 sky130_ef_ip__rdac3v_8bit_0/Vhigh ct2_switch_array_13/switch_array_2_0/channel1_in_to_out[1]
+ ct2_switch_array_13/switch_array_2_0/channel1_in_to_out[0] gpio_noesd[3] vdda1 vssa1
+ ct2_switch_array_13/switch_array_2_0/channel0_in_to_out[1] ct2_switch_array_13/switch_array_2_0/channel0_in_to_out[0]
+ sky130_ef_ip__rheostat_8bit_0/Vhigh vssd1 ct2_switch_array
Xsky130_ef_ip__cdac3v_12bit_0 sky130_ef_ip__cdac3v_12bit_0/SELD2 sky130_ef_ip__cdac3v_12bit_0/SELD3
+ sky130_ef_ip__cdac3v_12bit_0/SELD4 sky130_ef_ip__cdac3v_12bit_0/SELD5 sky130_ef_ip__cdac3v_12bit_0/SELD6
+ sky130_ef_ip__cdac3v_12bit_0/SELD7 sky130_ef_ip__cdac3v_12bit_0/SELD8 sky130_ef_ip__cdac3v_12bit_0/SELD9
+ io_analog[7] vccd2 sky130_ef_ip__cdac3v_12bit_0/OUT sky130_ef_ip__cdac3v_12bit_0/RST
+ sky130_ef_ip__cdac3v_12bit_0/SELD10 sky130_ef_ip__cdac3v_12bit_0/SELD11 sky130_ef_ip__cdac3v_12bit_0/OUTNC
+ sky130_ef_ip__cdac3v_12bit_0/SELD0 sky130_ef_ip__cdac3v_12bit_0/SELD1 sky130_ef_ip__cdac3v_12bit_0/VL
+ sky130_ef_ip__cdac3v_12bit_0/VH vssd2 vssa2 sky130_ef_ip__cdac3v_12bit
Xsky130_ef_ip__rdac3v_8bit_0 sky130_ef_ip__rdac3v_8bit_0/b0 sky130_ef_ip__rdac3v_8bit_0/b1
+ sky130_ef_ip__rdac3v_8bit_0/b2 sky130_ef_ip__rdac3v_8bit_0/b3 sky130_ef_ip__rdac3v_8bit_0/b4
+ sky130_ef_ip__rdac3v_8bit_0/b5 sky130_ef_ip__rdac3v_8bit_0/b6 sky130_ef_ip__rdac3v_8bit_0/b7
+ sky130_ef_ip__rdac3v_8bit_0/out io_analog[0] sky130_ef_ip__rdac3v_8bit_0/ena vccd1
+ sky130_ef_ip__rdac3v_8bit_0/Vhigh sky130_ef_ip__rdac3v_8bit_0/Vlow vssa1 vssd1 sky130_ef_ip__rdac3v_8bit
Xct2_switch_array_14 vccd1 sky130_ef_ip__samplehold_0/in ct2_switch_array_14/switch_array_2_0/channel1_in_to_out[1]
+ la_data_in[118] ct2_switch_array_14/switch_array_2_0/channel1_out vdda1 vssa1 ct2_switch_array_14/switch_array_2_0/channel0_in_to_out[1]
+ la_data_in[119] sky130_sw_ip__bgrref_por_0/porb_h[1] vssd1 ct2_switch_array
Xct2_switch_array_15 vccd1 sky130_icrg_ip__ulpcomp2_0/vinp ct2_switch_array_15/switch_array_2_0/channel1_in_to_out[1]
+ la_data_in[120] gpio_noesd[4] vdda1 vssa1 ct2_switch_array_15/switch_array_2_0/channel0_in_to_out[1]
+ ct2_switch_array_15/switch_array_2_0/channel0_in_to_out[0] sky130_aa_ip__programmable_pll_0/LF_OFFCHIP
+ vssd1 ct2_switch_array
Xsky130_ef_ip__rc_osc_500k_1 io_analog[4] vccd1 sky130_ef_ip__rc_osc_500k_1/ena io_out[13]
+ vssd1 vssa1 sky130_ef_ip__rc_osc_500k
R0 m3_800_463198# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R1 m3_800_333532# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R2 vssd1 m3_584112_456428# sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R3 m3_800_506420# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R4 gpio_analog[17] bias_reference_voltage sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
R5 vssd1 io_oeb[7] sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R6 vssd1 io_oeb[13] sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R7 m3_800_247288# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R8 sky130_ef_ip__rdac3v_8bit_0/Vhigh m3_583600_16528# sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R9 sky130_ef_ip__rdac3v_8bit_0/Vlow m3_583898_21256# sky130_fd_pr__res_generic_m3 w=0.56 l=0.63
R10 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R11 io_oeb[17] vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R12 m3_800_419976# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R13 m3_800_290310# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R14 sky130_ef_ip__rheostat_8bit_0/Vhigh m3_583894_47714# sky130_fd_pr__res_generic_m3 w=0.56 l=0.61
R15 sky130_ef_ip__rheostat_8bit_0/Vlow m3_584180_92372# sky130_fd_pr__res_generic_m3 w=0.56 l=0.52
R16 vssd1 m3_584000_412006# sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
R17 m3_800_119666# vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
R18 vssd1 io_oeb[8] sky130_fd_pr__res_generic_m3 w=0.56 l=0.56
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ io_analog[4]_uq0 io_analog[4]_uq1 io_analog[4]_uq2 io_analog[4]_uq3 io_analog[4]_uq4
+ io_analog[5]_uq0 io_analog[5]_uq1 io_analog[5]_uq2 io_analog[5]_uq3 io_analog[5]_uq4
+ io_analog[6]_uq0 io_analog[6]_uq1 io_analog[6]_uq2 io_analog[6]_uq3 io_analog[6]_uq4
+ vssa1 vssd2 vssd1 vssa2
Xchipalooza_testchip_2_0 gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17]
+ gpio_analog[1] gpio_analog[5] gpio_analog[6] gpio_analog[8] gpio_analog[9] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[7] io_analog[0] io_analog[10] io_analog[1]
+ io_analog[2] io_analog[3] io_analog[4]_uq3 io_analog[7] io_analog[8] io_analog[9]
+ io_analog[5]_uq4 io_analog[6]_uq4 io_oeb[0] io_oeb[12] io_oeb[13] io_oeb[17] io_oeb[1]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6]
+ io_oeb[7] io_oeb[8] io_out[0] io_out[12] io_out[13] io_out[17] io_out[1] io_out[23]
+ io_out[24] io_out[25] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[120] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[11] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] vccd1 vccd2 vdda1 vdda2 la_data_in[106] la_data_in[101] wbs_dat_i[6]
+ la_data_in[52] la_oenb[0] io_in[23] io_oeb[15] la_data_in[104] la_data_in[95] la_oenb[34]
+ wbs_dat_i[26] la_data_in[108] la_data_in[42] la_oenb[117] gpio_noesd[15] la_data_in[59]
+ wbs_dat_o[20] io_in_3v3[7] wbs_dat_o[12] gpio_analog[7] la_data_in[48] la_oenb[14]
+ io_in[14] gpio_noesd[9] wbs_dat_o[4] wbs_dat_o[7] wbs_sel_i[0] gpio_noesd[1] la_oenb[109]
+ la_data_in[78] la_oenb[98] wbs_dat_o[27] wbs_dat_i[4] la_data_in[115] io_in_3v3[15]
+ io_oeb[14] la_data_in[47] la_data_in[26] io_in_3v3[1] la_data_in[33] wbs_adr_i[22]
+ la_oenb[100] la_oenb[110] io_in[6] wbs_adr_i[14] la_data_in[40] io_analog[4]_uq2
+ la_data_in[12] gpio_analog[2] wbs_dat_o[18] la_oenb[85] io_oeb[10] wbs_we_i la_data_in[31]
+ la_oenb[74] wbs_dat_o[13] io_in_3v3[6] io_analog[6]_uq1 la_oenb[127] la_oenb[5]
+ io_in[20] io_in_3v3[26] la_oenb[123] la_data_in[17] la_data_in[65] la_oenb[102]
+ la_data_in[2] la_data_in[122] wbs_adr_i[20] la_oenb[19] la_data_in[57] wbs_adr_i[12]
+ la_data_in[41] io_in[13] la_data_in[93] wbs_dat_o[5] la_data_in[43] la_oenb[105]
+ wbs_adr_i[18] la_oenb[72] wbs_cyc_i wbs_dat_o[11] la_data_in[34] io_clamp_high[0]
+ wbs_dat_o[25] la_data_in[39] la_data_in[8] io_in_3v3[11] gpio_noesd[14] wbs_dat_o[31]
+ io_out[16] la_data_in[100] la_oenb[10] la_data_in[123] la_data_in[35] la_oenb[116]
+ io_in[2] la_oenb[83] la_data_in[110] io_in[21] la_data_in[50] wbs_sel_i[3] la_oenb[89]
+ la_data_in[91] wbs_adr_i[5] wbs_adr_i[16] io_in[18] la_oenb[20] wbs_dat_o[9] la_oenb[15]
+ gpio_analog[3] wbs_adr_i[25] io_analog[5]_uq1 io_out[22] gpio_noesd[10] user_irq[2]
+ la_data_in[28] wbs_dat_o[29] gpio_noesd[13] io_in_3v3[19] la_oenb[4] la_oenb[28]
+ io_oeb[18] la_oenb[111] la_data_in[121] la_oenb[21] wbs_dat_o[24] wbs_adr_i[24]
+ wbs_adr_i[19] wbs_adr_i[11] la_oenb[120] la_data_in[103] la_data_in[13] wbs_dat_i[2]
+ io_in[5] la_oenb[87] la_data_in[37] wbs_dat_i[3] la_oenb[6] io_oeb[26] io_in[10]
+ la_data_in[94] la_oenb[76] io_in[24] wbs_adr_i[31] la_oenb[46] la_oenb[3] la_oenb[71]
+ gpio_noesd[6] wbs_adr_i[3] io_out[14] la_oenb[30] la_data_in[125] io_in[4] wbs_dat_i[23]
+ la_data_in[46] wbs_adr_i[17] wb_clk_i io_analog[4] io_in_3v3[12] la_data_in[18]
+ wbs_sel_i[1] wbs_adr_i[23] io_analog[6]_uq2 la_oenb[63] la_oenb[80] user_irq[0]
+ la_oenb[69] wbs_adr_i[29] io_analog[6]_uq0 io_out[20] la_data_in[9] la_oenb[75]
+ io_clamp_low[2] gpio_noesd[11] user_clock2 la_oenb[11] wbs_adr_i[9] la_oenb[118]
+ io_oeb[11] wbs_dat_i[21] la_oenb[88] wbs_adr_i[15] io_out[18] wbs_adr_i[7] la_oenb[114]
+ wbs_adr_i[21] la_oenb[113] la_oenb[61] la_oenb[25] wbs_dat_o[1] la_oenb[86] la_data_in[23]
+ la_data_out[126] la_oenb[67] wbs_adr_i[27] la_data_in[96] io_in_3v3[16] io_in_3v3[8]
+ la_oenb[37] io_clamp_high[2] io_oeb[16] io_oeb[9] wbs_dat_i[16] wbs_dat_o[26] la_data_in[0]
+ io_out[10] gpio_noesd[16] wbs_dat_i[8] io_in[15] wbs_dat_o[2] wbs_adr_i[13] io_out[15]
+ wbs_dat_i[14] la_oenb[78] io_in[9] la_data_in[126] io_in[11] la_data_in[69] wbs_adr_i[8]
+ gpio_noesd[17] io_in_3v3[22] la_oenb[59] la_data_in[102] la_oenb[7] io_analog[5]_uq2
+ la_oenb[84] la_oenb[48] la_oenb[54] la_oenb[73] la_oenb[65] wbs_adr_i[28] la_oenb[43]
+ io_analog[5]_uq0 la_oenb[16] la_oenb[60] wbs_dat_i[22] la_data_in[124] wbs_dat_i[0]
+ la_oenb[94] la_data_in[32] la_data_in[80] io_clamp_low[1] la_oenb[122] io_in_3v3[18]
+ la_data_in[116] la_data_in[109] io_in[0] la_oenb[35] wbs_adr_i[1] la_data_in[86]
+ wbs_adr_i[0] la_data_in[1] gpio_noesd[0] la_data_in[75] la_oenb[125] la_oenb[90]
+ wbs_adr_i[6] la_data_in[105] gpio_noesd[12] la_oenb[68] la_data_in[19] la_data_in[112]
+ io_in_3v3[13] la_oenb[82] la_oenb[91] la_data_in[21] la_oenb[52] wbs_adr_i[26] la_oenb[95]
+ la_data_in[29] la_oenb[41] la_oenb[99] la_data_out[117] wbs_dat_i[20] la_oenb[26]
+ io_out[21] la_oenb[47] wbs_dat_i[12] la_data_in[67] la_oenb[2] io_in_3v3[23] la_data_in[84]
+ la_oenb[31] wbs_dat_o[0] la_data_in[10] io_analog[4]_uq1 la_oenb[97] la_oenb[108]
+ io_in[26] la_data_in[73] la_oenb[77] la_data_in[45] la_data_out[0] la_oenb[66] io_in_3v3[9]
+ la_data_in[5] io_in[7] io_analog[6] la_data_in[53] la_oenb[58] io_in_3v3[14] la_oenb[50]
+ la_oenb[39] la_oenb[96] la_oenb[64] gpio_noesd[5] wbs_dat_i[18] wbs_dat_o[19] la_oenb[45]
+ la_data_in[15] wbs_stb_i la_oenb[106] io_oeb[22] gpio_noesd[8] wbs_dat_i[10] wbs_dat_i[13]
+ wbs_dat_i[24] la_data_in[30] io_in[19] la_oenb[33] wbs_dat_i[27] la_oenb[40] io_in[1]
+ wbs_adr_i[4] io_oeb[20] la_oenb[12] la_data_in[90] la_data_in[27] la_data_in[111]
+ la_data_in[4] wbs_dat_i[19] la_data_in[71] wbs_adr_i[10] io_in_3v3[4] la_data_in[66]
+ wbs_dat_i[25] io_oeb[19] la_oenb[24] la_oenb[56] io_in_3v3[10] la_oenb[70] la_oenb[107]
+ wbs_adr_i[30] la_oenb[101] la_oenb[126] la_data_in[6] la_oenb[62] wbs_dat_i[5] la_oenb[17]
+ io_out[19] wbs_dat_o[17] la_data_in[82] wbs_dat_i[11] la_data_in[25] la_oenb[115]
+ io_in[12] io_out[9] la_oenb[103] la_data_in[88] la_data_in[92] wbs_dat_o[3] la_data_in[58]
+ la_data_in[77] la_oenb[81] wbs_dat_i[31] io_out[11] la_data_in[83] la_data_out[24]
+ la_data_in[14] la_data_in[54] la_oenb[29] la_data_in[72] la_data_in[64] la_data_out[127]
+ io_analog[5] la_oenb[57] io_in_3v3[25] la_oenb[22] la_oenb[8] la_data_in[98] io_in[17]
+ la_data_out[119] wbs_ack_o la_oenb[49] la_oenb[112] la_data_in[24] io_clamp_low[0]
+ la_oenb[38] wbs_dat_i[17] wbs_dat_i[9] wb_rst_i la_oenb[23] la_data_in[114] la_data_in[89]
+ wbs_adr_i[2] la_data_in[56] la_oenb[79] wbs_dat_i[29] la_data_in[11] io_in_3v3[21]
+ la_oenb[13] la_data_in[81] user_irq[1] la_oenb[32] io_oeb[21] la_data_in[70] io_in[25]
+ io_analog[4]_uq4 la_data_in[51] io_in[8] wbs_dat_o[23] la_data_in[107] la_oenb[27]
+ la_oenb[55] wbs_dat_o[15] io_in_3v3[2] la_oenb[44] io_in_3v3[3] la_oenb[92] io_analog[6]_uq3
+ io_in[22] wbs_dat_o[10] la_oenb[36] wbs_dat_o[21] la_data_in[3] io_in[16] wbs_dat_i[15]
+ la_oenb[93] la_oenb[42] la_data_in[113] wbs_dat_o[30] la_oenb[1] la_data_in[62]
+ la_data_in[76] io_in_3v3[17] io_analog[4]_uq0 io_in[3] la_data_in[79] la_data_in[49]
+ la_data_in[68] wbs_dat_i[30] la_data_in[99] la_data_in[44] io_out[26] la_data_out[120]
+ la_data_in[38] io_in_3v3[24] la_data_in[127] wbs_dat_o[16] la_oenb[53] la_data_in[22]
+ wbs_dat_i[7] la_oenb[121] la_data_in[7] wbs_dat_o[8] wbs_dat_o[22] la_data_in[87]
+ wbs_sel_i[2] io_clamp_high[1] io_in_3v3[5] la_data_in[16] wbs_dat_o[28] la_data_in[60]
+ w_532863_486748# la_data_in[63] la_data_in[74] la_oenb[18] io_in_3v3[0] la_oenb[124]
+ la_data_in[55] gpio_analog[4] wbs_dat_i[28] la_data_in[20] la_data_out[118] la_oenb[104]
+ la_data_in[36] io_in_3v3[20] la_oenb[119] la_data_in[61] wbs_dat_o[14] la_oenb[51]
+ la_oenb[9] vssd1 vssd2 wbs_dat_o[6] la_data_in[97] gpio_analog[8] vssa2 vssa1 la_data_in[85]
+ io_analog[5]_uq3 wbs_dat_i[1] chipalooza_testchip_2
.ends

