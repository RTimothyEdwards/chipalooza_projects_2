magic
tech sky130A
magscale 1 2
timestamp 1726424352
<< isosubstrate >>
rect 800 649262 286990 704800
rect 800 602768 170886 649262
rect 800 593672 23894 602768
rect 68592 593672 170886 602768
rect 800 574516 23826 593672
rect 73604 574516 170886 593672
rect 800 565418 23894 574516
rect 67046 574016 170886 574516
rect 246186 645696 286990 649262
rect 246186 638532 247860 645696
rect 264682 638532 286990 645696
rect 246186 574016 286990 638532
rect 67046 565418 286990 574016
rect 800 559252 286990 565418
rect 800 523928 170874 559252
rect 800 511962 3562 523928
rect 9554 516322 170874 523928
rect 9554 511962 33612 516322
rect 800 497388 33612 511962
rect 800 492344 35896 497388
rect 51126 492344 170874 516322
rect 800 484006 170874 492344
rect 246156 555704 286990 559252
rect 246156 548548 247878 555704
rect 264686 548548 286990 555704
rect 246156 484006 286990 548548
rect 800 480808 286990 484006
rect 800 468842 3562 480808
rect 9592 469242 286990 480808
rect 9592 468842 170882 469242
rect 800 437584 170882 468842
rect 800 425618 3562 437584
rect 9574 433426 170882 437584
rect 9574 425618 39254 433426
rect 52414 426808 170882 433426
rect 800 413468 39254 425618
rect 49484 424166 170882 426808
rect 52426 413468 170882 424166
rect 800 394292 170882 413468
rect 800 382326 3528 394292
rect 9564 394008 170882 394292
rect 246182 465714 286990 469242
rect 246182 458550 247860 465714
rect 264688 458550 286990 465714
rect 246182 394008 286990 458550
rect 9564 382326 286990 394008
rect 800 379244 286990 382326
rect 800 350762 170902 379244
rect 800 338796 3494 350762
rect 9582 340440 170902 350762
rect 9582 338796 24996 340440
rect 800 327542 24996 338796
rect 35724 336394 170902 340440
rect 36518 327542 170902 336394
rect 800 307846 170902 327542
rect 800 295880 3562 307846
rect 9554 304002 170902 307846
rect 246174 375710 286990 379244
rect 246174 368538 247864 375710
rect 264690 368538 286990 375710
rect 246174 304002 286990 368538
rect 9554 295880 286990 304002
rect 800 289254 286990 295880
rect 800 274518 170880 289254
rect 800 272642 24830 274518
rect 800 268614 30198 272642
rect 61422 272618 170880 274518
rect 56364 268624 170880 272618
rect 800 265618 24830 268614
rect 61422 265618 170880 268624
rect 800 264760 30188 265618
rect 800 252794 3494 264760
rect 9574 261624 30188 264760
rect 56308 261624 170880 265618
rect 9574 258604 24980 261624
rect 9574 254610 30188 258604
rect 61422 258594 170880 261624
rect 9574 252794 25048 254610
rect 56318 254600 170880 258594
rect 800 251626 25048 252794
rect 800 251352 30098 251626
rect 61422 251614 170880 254600
rect 800 247850 30144 251352
rect 800 247610 30098 247850
rect 56374 247620 170880 251614
rect 800 244602 24992 247610
rect 61422 244624 170880 247620
rect 800 244314 30142 244602
rect 800 240776 30144 244314
rect 800 240630 30142 240776
rect 56352 240630 170880 244624
rect 800 237612 25038 240630
rect 61422 237636 170880 240630
rect 800 233606 30176 237612
rect 56352 233618 170880 237636
rect 800 230600 25004 233606
rect 61422 230612 170880 233618
rect 800 226616 30176 230600
rect 800 224650 25038 226616
rect 56308 226594 170880 230612
rect 61422 224650 170880 226594
rect 800 214012 170880 224650
rect 246176 285712 286990 289254
rect 246176 278532 247850 285712
rect 264684 278532 286990 285712
rect 246176 214012 286990 278532
rect 800 199234 286990 214012
rect 800 137316 170880 199234
rect 800 125350 4008 137316
rect 10154 135214 170880 137316
rect 10154 131168 30558 135214
rect 42054 131324 170880 135214
rect 10154 125350 30592 131168
rect 39926 129024 170880 131324
rect 800 125208 30592 125350
rect 42230 125208 170880 129024
rect 800 124014 170880 125208
rect 246178 195706 286990 199234
rect 246178 188532 247860 195706
rect 264692 188532 286990 195706
rect 246178 124014 286990 188532
rect 800 109252 286990 124014
rect 800 94128 170888 109252
rect 800 82162 4008 94128
rect 10116 82162 170888 94128
rect 800 73686 170888 82162
rect 800 50644 30166 73686
rect 800 38678 4044 50644
rect 10146 43988 30166 50644
rect 40740 43988 170888 73686
rect 10146 38678 170888 43988
rect 800 34020 170888 38678
rect 246172 105696 286990 109252
rect 246172 98536 247842 105696
rect 264664 98536 286990 105696
rect 246172 34020 286990 98536
rect 800 800 286990 34020
rect 296274 649224 584800 704800
rect 296274 645702 340588 649224
rect 296274 638542 322086 645702
rect 338916 638542 340588 645702
rect 296274 574012 340588 638542
rect 415890 617042 584800 649224
rect 415890 612192 545950 617042
rect 559260 612364 584800 617042
rect 415890 605408 545986 612192
rect 556652 610288 584800 612364
rect 559152 605408 584800 610288
rect 415890 598548 584800 605408
rect 415890 586408 574674 598548
rect 581230 586408 584800 598548
rect 415890 574012 584800 586408
rect 296274 559230 584800 574012
rect 296274 555702 340592 559230
rect 296274 548546 322096 555702
rect 338924 548546 340592 555702
rect 296274 484020 340592 548546
rect 415900 523914 584800 559230
rect 415900 519678 537218 523914
rect 548188 519678 584800 523914
rect 415900 519334 584800 519678
rect 415900 513728 533764 519334
rect 536398 518648 584800 519334
rect 536398 514430 537226 518648
rect 548214 517830 584800 518648
rect 548214 514430 574918 517830
rect 536398 513728 574918 514430
rect 415900 505690 574918 513728
rect 581302 505690 584800 517830
rect 415900 501436 584800 505690
rect 415900 489420 574906 501436
rect 415900 487054 533224 489420
rect 537996 489296 574906 489420
rect 581374 489296 584800 501436
rect 537996 487054 584800 489296
rect 415900 484970 584800 487054
rect 415900 484020 574944 484970
rect 296274 472830 574944 484020
rect 581266 472830 584800 484970
rect 296274 469234 584800 472830
rect 296274 465716 340584 469234
rect 296274 458548 322090 465716
rect 338916 458548 340584 465716
rect 296274 394018 340584 458548
rect 415880 394018 584800 469234
rect 296274 379250 584800 394018
rect 296274 375706 340592 379250
rect 296274 368532 322092 375706
rect 338910 368532 340592 375706
rect 296274 304010 340592 368532
rect 415902 323436 584800 379250
rect 415902 311590 574906 323436
rect 581132 311590 584800 323436
rect 415902 304010 584800 311590
rect 296274 289228 584800 304010
rect 296274 285712 340602 289228
rect 296274 278540 322084 285712
rect 338922 278540 340602 285712
rect 296274 214030 340602 278540
rect 415902 284094 584800 289228
rect 415902 272248 574932 284094
rect 581132 272248 584800 284094
rect 415902 260230 584800 272248
rect 415902 253134 527695 260230
rect 541403 253134 584800 260230
rect 415902 214030 584800 253134
rect 296274 199236 584800 214030
rect 296274 195702 340588 199236
rect 296274 188538 322092 195702
rect 338916 188538 340588 195702
rect 296274 124012 340588 188538
rect 415874 181204 584800 199236
rect 415874 160034 534250 181204
rect 550970 160034 584800 181204
rect 415874 124012 584800 160034
rect 296274 109274 584800 124012
rect 296274 105696 340616 109274
rect 296274 98536 322088 105696
rect 338914 98536 340616 105696
rect 296274 34000 340616 98536
rect 415896 83024 584800 109274
rect 415896 62068 535616 83024
rect 552282 80162 584800 83024
rect 552282 69200 553252 80162
rect 557468 69200 584800 80162
rect 552282 62068 584800 69200
rect 415896 34000 584800 62068
rect 296274 800 584800 34000
<< locali >>
rect 466566 388495 466798 388631
rect 467018 386128 467320 386264
rect 467262 385111 467680 385247
rect 461455 382166 461615 382200
rect 486342 380902 486440 380966
rect 477002 379426 477054 379496
rect 461599 377587 462997 377841
rect 461657 377189 462867 377479
rect 461904 376009 462924 376421
rect 461941 374677 462789 375111
rect 559447 373108 561334 376077
rect 577998 368301 580967 371074
rect 448496 368180 449236 368196
rect 448496 367479 448509 368180
rect 449223 367479 449236 368180
rect 519860 367938 520094 367944
rect 519860 367870 519866 367938
rect 519934 367870 520094 367938
rect 519860 367864 520094 367870
rect 448496 367464 449236 367479
rect 448991 364753 449547 364883
rect 477802 352726 478234 352862
rect 477852 352527 478534 352663
rect 477768 352294 478884 352430
rect 477734 352039 479216 352175
rect 477768 351753 479600 351889
rect 477868 351454 479900 351590
rect 477734 351084 480282 351220
rect 477734 350840 480664 350976
rect 449761 347585 450162 347803
rect 449334 329928 449792 330107
rect 449370 317337 449574 317473
<< viali >>
rect 466798 388495 466934 388631
rect 466938 387792 467074 387928
rect 467320 386128 467456 386264
rect 467680 385111 467816 385247
rect 478342 382470 478416 382544
rect 461421 382166 461455 382200
rect 477002 379374 477054 379426
rect 461345 377587 461599 377841
rect 461367 377189 461657 377479
rect 461492 376009 461904 376421
rect 461507 374677 461941 375111
rect 556478 373108 559447 376077
rect 448467 371062 449133 371715
rect 448509 367479 449223 368180
rect 519866 367870 519934 367938
rect 577998 365332 580967 368301
rect 448861 364753 448991 364883
rect 478234 352726 478370 352862
rect 478534 352527 478670 352663
rect 478884 352294 479020 352430
rect 479216 352039 479352 352175
rect 479600 351753 479736 351889
rect 479900 351454 480036 351590
rect 480282 351084 480418 351220
rect 480664 350840 480800 350976
rect 449543 347585 449761 347803
rect 457398 336135 457534 336271
rect 457082 335936 457218 336072
rect 456768 335703 456904 335839
rect 456452 335448 456588 335584
rect 449155 329928 449334 330107
rect 451918 318024 452054 318160
rect 450034 317825 450170 317961
rect 449672 317592 449808 317728
rect 449234 317337 449370 317473
<< metal1 >>
rect 265195 657031 265674 657037
rect 246223 655231 247829 655237
rect 246223 647742 247829 653625
rect 265195 648452 265674 656552
rect 321112 657031 321591 657037
rect 321112 648931 321591 656552
rect 338957 655231 340563 655237
rect 338957 649354 340563 653625
rect 338957 649320 340644 649354
rect 338957 649280 340599 649320
rect 338957 649254 340644 649280
rect 321112 648930 321596 648931
rect 321117 648904 321596 648930
rect 338957 647712 340599 649254
rect 338962 647592 340568 647712
rect 340573 647592 340599 647712
rect 558396 612276 561641 612654
rect 558396 609925 560291 610303
rect 560669 609925 560675 610303
rect 561263 610291 561641 612276
rect 561263 609907 561641 609913
rect 72086 597575 72802 597643
rect 72870 597575 72876 597643
rect 72078 595947 72744 596015
rect 72812 595947 72818 596015
rect 72050 593643 76475 593764
rect 76596 593643 76602 593764
rect 265195 567031 265674 567037
rect 246223 565231 247829 565237
rect 246223 559354 247829 563625
rect 246086 559320 247829 559354
rect 246192 559280 246218 559320
rect 246086 559254 246218 559280
rect 246192 557712 246218 559254
rect 246223 557712 247829 559320
rect 265195 558930 265674 566552
rect 321112 567031 321591 567037
rect 321112 558931 321591 566552
rect 338957 565231 340563 565237
rect 338957 559354 340563 563625
rect 338957 559320 340644 559354
rect 338957 559280 340599 559320
rect 338957 559254 340644 559280
rect 321112 558930 321596 558931
rect 321117 558904 321596 558930
rect 338957 557712 340599 559254
rect 338962 557592 340568 557712
rect 340573 557592 340599 557712
rect 532580 522710 532586 522794
rect 532670 522710 534138 522794
rect 532504 520206 532510 520290
rect 532594 520206 534086 520290
rect 530211 501689 530297 501695
rect 530211 481564 530297 501603
rect 530691 501161 530697 501247
rect 530783 501161 530789 501247
rect 530697 483196 530783 501161
rect 541778 488174 544533 488260
rect 544619 488174 544625 488260
rect 530697 483110 532781 483196
rect 542128 481586 542134 481594
rect 530211 481478 532914 481564
rect 541590 481550 542134 481586
rect 542128 481542 542134 481550
rect 542186 481586 542192 481594
rect 542186 481550 542214 481586
rect 542186 481542 542192 481550
rect 541952 480668 542004 480674
rect 541590 480624 541952 480660
rect 542004 480624 542032 480660
rect 541952 480610 542004 480616
rect 265195 477031 265674 477037
rect 246223 475231 247829 475237
rect 246223 469354 247829 473625
rect 246086 469320 247829 469354
rect 246192 469280 246218 469320
rect 246086 469254 246218 469280
rect 246192 467712 246218 469254
rect 246223 467712 247829 469320
rect 265195 468930 265674 476552
rect 321112 477031 321591 477037
rect 321112 468931 321591 476552
rect 338957 475231 340563 475237
rect 338957 469354 340563 473625
rect 338957 469320 340644 469354
rect 338957 469280 340599 469320
rect 338957 469254 340644 469280
rect 321112 468930 321596 468931
rect 321117 468904 321596 468930
rect 338957 467712 340599 469254
rect 338962 467592 340568 467712
rect 340573 467592 340599 467712
rect 52496 426798 52785 426872
rect 52859 426798 53198 426872
rect 52504 426508 52877 426582
rect 52951 426508 53206 426582
rect 52320 426023 52894 426223
rect 53094 426023 53100 426223
rect 52484 425596 53035 425670
rect 53109 425596 53186 425670
rect 52478 425314 53043 425388
rect 53117 425314 53180 425388
rect 52474 425042 53035 425116
rect 53109 425042 53176 425116
rect 52321 424701 53034 424901
rect 53234 424701 53240 424901
rect 52321 424396 53034 424596
rect 53234 424396 53240 424596
rect 34440 423301 34446 423501
rect 34646 423301 39401 423501
rect 33744 423001 33750 423201
rect 33950 423001 39401 423201
rect 33034 422901 33234 422907
rect 33234 422701 39401 422901
rect 33034 422695 33234 422701
rect 32362 422601 32562 422607
rect 32562 422401 39401 422601
rect 32362 422395 32562 422401
rect 37902 422101 37908 422301
rect 38108 422101 39404 422301
rect 466792 388631 466940 388643
rect 466792 388495 466798 388631
rect 466934 388495 467308 388631
rect 467444 388495 467450 388631
rect 466792 388483 466940 388495
rect 466924 387928 467088 387934
rect 466924 387792 466938 387928
rect 467074 387792 467298 387928
rect 467434 387792 467440 387928
rect 466924 387786 467088 387792
rect 265195 387031 265674 387037
rect 246223 385231 247829 385237
rect 246223 379354 247829 383625
rect 246086 379320 247829 379354
rect 246192 379280 246218 379320
rect 246086 379254 246218 379280
rect 246192 377712 246218 379254
rect 246223 377712 247829 379320
rect 265195 378930 265674 386552
rect 321112 387031 321591 387037
rect 321112 378931 321591 386552
rect 467314 386264 467462 386276
rect 467314 386128 467320 386264
rect 467456 386128 467912 386264
rect 468048 386128 468054 386264
rect 467314 386116 467462 386128
rect 467674 385247 467822 385259
rect 338957 385231 340563 385237
rect 467674 385111 467680 385247
rect 467816 385111 468168 385247
rect 468304 385111 468310 385247
rect 467674 385099 467822 385111
rect 338957 379354 340563 383625
rect 478342 383269 478416 383275
rect 478342 382564 478416 383195
rect 478336 382544 478422 382564
rect 478336 382470 478342 382544
rect 478416 382470 478422 382544
rect 478336 382458 478422 382470
rect 461118 382209 461170 382215
rect 461415 382200 461461 382212
rect 461170 382166 461421 382200
rect 461455 382166 461461 382200
rect 461118 382151 461170 382157
rect 461415 382154 461461 382166
rect 464333 381270 464469 381630
rect 458190 381134 458196 381270
rect 458332 381134 464469 381270
rect 486342 380959 486440 380966
rect 486342 380907 486382 380959
rect 486434 380907 486440 380959
rect 486342 380902 486440 380907
rect 476990 379426 477066 379432
rect 476990 379374 477002 379426
rect 477054 379374 477066 379426
rect 476990 379368 477066 379374
rect 338957 379320 340644 379354
rect 338957 379280 340599 379320
rect 338957 379254 340644 379280
rect 321112 378930 321596 378931
rect 321117 378904 321596 378930
rect 338957 377712 340599 379254
rect 477002 379226 477054 379368
rect 477002 379168 477054 379174
rect 486574 378502 488527 378596
rect 488621 378502 488627 378596
rect 480832 378274 483683 378368
rect 483777 378274 483783 378368
rect 485662 377992 487669 378086
rect 487763 377992 487769 378086
rect 461339 377841 461605 377853
rect 338962 377592 340568 377712
rect 340573 377592 340599 377712
rect 459329 377587 459335 377841
rect 459589 377587 461345 377841
rect 461599 377587 461605 377841
rect 461339 377575 461605 377587
rect 461361 377479 461663 377491
rect 459525 377189 459531 377479
rect 459821 377189 461367 377479
rect 461657 377189 461663 377479
rect 461361 377177 461663 377189
rect 501381 377151 501711 377157
rect 461486 376421 461910 376433
rect 459778 376009 459784 376421
rect 460196 376009 461492 376421
rect 461904 376009 461910 376421
rect 501381 376131 501711 376821
rect 556472 376077 559453 376089
rect 461486 375997 461910 376009
rect 500454 375546 500534 375552
rect 518984 375546 519064 375552
rect 502386 375466 502392 375546
rect 502472 375466 518984 375546
rect 500454 375460 500534 375466
rect 518984 375460 519064 375466
rect 461501 375111 461947 375123
rect 459859 374677 459865 375111
rect 460299 374677 461507 375111
rect 461941 374677 461947 375111
rect 461501 374665 461947 374677
rect 502022 372934 502102 373364
rect 553596 373108 553602 376077
rect 559447 373108 559453 376077
rect 556472 373096 559453 373108
rect 520746 372934 520826 372940
rect 502022 372854 520746 372934
rect 520746 372848 520826 372854
rect 448461 371715 449139 371721
rect 442628 371062 442634 371715
rect 443287 371062 448467 371715
rect 449133 371062 450906 371715
rect 448461 371056 449139 371062
rect 577986 368301 580979 368307
rect 448496 368180 449236 368196
rect 441438 367479 441444 368180
rect 442145 367479 448509 368180
rect 449223 367479 449236 368180
rect 520840 367944 520920 367950
rect 519854 367938 520840 367944
rect 519854 367870 519866 367938
rect 519934 367870 520840 367938
rect 519854 367864 520840 367870
rect 520840 367858 520920 367864
rect 448496 367464 449236 367479
rect 577986 365332 577998 368301
rect 580967 365332 580979 368301
rect 577986 365326 580979 365332
rect 448855 364883 448997 364895
rect 439827 364753 439833 364883
rect 439963 364753 448861 364883
rect 448991 364753 448997 364883
rect 448855 364741 448997 364753
rect 577998 363733 580967 365326
rect 577998 360758 580967 360764
rect 478222 352862 478382 352868
rect 478222 352726 478234 352862
rect 478370 352726 478382 352862
rect 478222 352720 478382 352726
rect 439337 347803 439555 347809
rect 449537 347803 449767 347815
rect 439555 347585 449543 347803
rect 449761 347585 449767 347803
rect 439337 347579 439555 347585
rect 449537 347573 449767 347585
rect 478234 347302 478370 352720
rect 478528 352663 478676 352675
rect 478528 352527 478534 352663
rect 478670 352527 478676 352663
rect 478528 352515 478676 352527
rect 478534 347572 478670 352515
rect 478878 352430 479026 352442
rect 478878 352294 478884 352430
rect 479020 352294 479026 352430
rect 478878 352282 479026 352294
rect 478884 347842 479020 352282
rect 479204 352175 479364 352181
rect 479204 352039 479216 352175
rect 479352 352039 479364 352175
rect 479204 352033 479364 352039
rect 479216 348096 479352 352033
rect 479594 351889 479742 351901
rect 479594 351753 479600 351889
rect 479736 351753 479742 351889
rect 479594 351741 479742 351753
rect 479600 348366 479736 351741
rect 479894 351590 480042 351602
rect 479894 351454 479900 351590
rect 480036 351454 480042 351590
rect 479894 351442 480042 351454
rect 479900 348720 480036 351442
rect 480276 351220 480424 351232
rect 480276 351084 480282 351220
rect 480418 351084 480424 351220
rect 480276 351072 480424 351084
rect 480282 349058 480418 351072
rect 480658 350976 480806 350988
rect 480658 350840 480664 350976
rect 480800 350840 480806 350976
rect 480658 350828 480806 350840
rect 480664 349378 480800 350828
rect 480664 349242 483026 349378
rect 483162 349242 483168 349378
rect 480664 349220 480800 349242
rect 483044 349058 483180 349064
rect 480282 348922 483044 349058
rect 483044 348916 483180 348922
rect 479900 348584 483044 348720
rect 483180 348584 483186 348720
rect 483078 348366 483214 348372
rect 479600 348230 483078 348366
rect 483078 348224 483214 348230
rect 479216 347960 483094 348096
rect 483230 347960 483236 348096
rect 478884 347706 483128 347842
rect 483264 347706 483270 347842
rect 483178 347572 483314 347578
rect 478534 347436 483178 347572
rect 483178 347430 483314 347436
rect 483212 347302 483348 347308
rect 478234 347166 483212 347302
rect 483212 347160 483348 347166
rect 38117 340222 38169 340228
rect 38117 339956 38169 340170
rect 457392 336271 457540 336288
rect 457392 336135 457398 336271
rect 457534 336135 457540 336271
rect 457392 336120 457540 336135
rect 457076 336072 457224 336090
rect 457076 335936 457082 336072
rect 457218 335936 457224 336072
rect 457076 335920 457224 335936
rect 456762 335839 456910 335856
rect 456762 335703 456768 335839
rect 456904 335703 456910 335839
rect 456762 335690 456910 335703
rect 456446 335584 456594 335602
rect 456446 335448 456452 335584
rect 456588 335448 456594 335584
rect 456446 335434 456594 335448
rect 449149 330107 449340 330119
rect 438557 329928 438563 330107
rect 438742 329928 449155 330107
rect 449334 329928 449340 330107
rect 449149 329916 449340 329928
rect 451912 318160 452060 318178
rect 451912 318024 451918 318160
rect 452054 318024 452060 318160
rect 451912 318010 452060 318024
rect 450028 317961 450176 317980
rect 450028 317825 450034 317961
rect 450170 317825 450176 317961
rect 450028 317810 450176 317825
rect 449666 317728 449814 317748
rect 449666 317592 449672 317728
rect 449808 317592 449814 317728
rect 449666 317578 449814 317592
rect 449228 317473 449376 317496
rect 449228 317337 449234 317473
rect 449370 317337 449376 317473
rect 449228 317314 449376 317337
rect 449234 310732 449370 317314
rect 449672 311266 449808 317578
rect 450034 311702 450170 317810
rect 451918 312270 452054 318010
rect 456452 312838 456588 335434
rect 456768 313174 456904 335690
rect 457082 313542 457218 335920
rect 457398 314010 457534 336120
rect 457398 313970 519868 314010
rect 457398 313890 519754 313970
rect 519834 313890 519868 313970
rect 457398 313874 519868 313890
rect 457082 313516 519692 313542
rect 457082 313436 519594 313516
rect 519674 313436 519692 313516
rect 457082 313406 519692 313436
rect 456768 313164 519542 313174
rect 456768 313084 519434 313164
rect 519514 313084 519542 313164
rect 456768 313038 519542 313084
rect 456452 312776 519398 312838
rect 456452 312702 519274 312776
rect 519268 312696 519274 312702
rect 519354 312702 519398 312776
rect 519354 312696 519360 312702
rect 451918 312230 519188 312270
rect 451918 312150 519054 312230
rect 519134 312150 519188 312230
rect 451918 312134 519188 312150
rect 450034 311660 519020 311702
rect 450034 311580 518894 311660
rect 518974 311580 519020 311660
rect 450034 311566 519020 311580
rect 449672 311230 518836 311266
rect 449672 311150 518734 311230
rect 518814 311150 518836 311230
rect 449672 311130 518836 311150
rect 449234 310692 518692 310732
rect 449234 310612 518574 310692
rect 518654 310612 518692 310692
rect 449234 310596 518692 310612
rect 265195 297031 265674 297037
rect 246223 295231 247829 295237
rect 246223 289354 247829 293625
rect 246086 289320 247829 289354
rect 246192 289280 246218 289320
rect 246086 289254 246218 289280
rect 246192 287712 246218 289254
rect 246223 287712 247829 289320
rect 265195 288930 265674 296552
rect 321112 297031 321591 297037
rect 321112 288931 321591 296552
rect 338957 295231 340563 295237
rect 338957 289354 340563 293625
rect 338957 289320 340644 289354
rect 338957 289280 340599 289320
rect 338957 289254 340644 289280
rect 321112 288930 321596 288931
rect 321117 288904 321596 288930
rect 338957 287712 340599 289254
rect 338962 287592 340568 287712
rect 340573 287592 340599 287712
rect 265195 207031 265674 207037
rect 246223 205231 247829 205237
rect 246223 199354 247829 203625
rect 246086 199320 247829 199354
rect 246192 199280 246218 199320
rect 246086 199254 246218 199280
rect 246192 197712 246218 199254
rect 246223 197712 247829 199320
rect 265195 198930 265674 206552
rect 321112 207031 321591 207037
rect 321112 198931 321591 206552
rect 338957 205231 340563 205237
rect 338957 199354 340563 203625
rect 338957 199320 340644 199354
rect 338957 199280 340599 199320
rect 338957 199254 340644 199280
rect 321112 198930 321596 198931
rect 321117 198904 321596 198930
rect 338957 197712 340599 199254
rect 338962 197592 340568 197712
rect 340573 197592 340599 197712
rect 551624 170290 552198 170461
rect 552369 170290 552375 170461
rect 535443 152725 535501 154707
rect 535443 152661 535501 152667
rect 537071 152493 537129 154697
rect 537071 152429 537129 152435
rect 538699 152343 538757 154693
rect 538699 152279 538757 152285
rect 540327 152179 540385 154679
rect 540327 152115 540385 152121
rect 541955 152025 542013 154674
rect 541955 151961 542013 151967
rect 543583 151787 543641 154675
rect 543583 151723 543641 151729
rect 545211 151633 545269 154675
rect 545211 151569 545269 151575
rect 546839 151475 546897 154675
rect 546839 151411 546897 151417
rect 41424 131168 43657 131546
rect 44035 131168 44041 131546
rect 41424 128787 43661 129165
rect 44039 128787 44045 129165
rect 265195 117031 265674 117037
rect 246223 115231 247829 115237
rect 246223 109354 247829 113625
rect 246086 109320 247829 109354
rect 246192 109280 246218 109320
rect 246086 109254 246218 109280
rect 246192 107712 246218 109254
rect 246223 107712 247829 109320
rect 265195 108930 265674 116552
rect 321112 117031 321591 117037
rect 321112 108930 321591 116552
rect 338957 115231 340563 115237
rect 338957 109354 340563 113625
rect 338957 109320 340700 109354
rect 338957 107712 340563 109320
rect 340568 109280 340594 109320
rect 340568 109254 340700 109280
rect 340568 107712 340594 109254
rect 40010 59508 40182 59528
rect 40010 58154 40028 59508
rect 40164 58154 40182 59508
rect 40010 58138 40182 58154
rect 536995 56509 537053 56515
rect 536995 56445 537053 56451
rect 538623 56385 538681 56523
rect 540251 56407 540309 56541
rect 540251 56343 540309 56349
rect 541879 56389 541937 56535
rect 538623 56321 538681 56327
rect 541879 56325 541937 56331
rect 543507 56325 543565 56523
rect 543507 56261 543565 56267
rect 545135 56197 545193 56567
rect 546763 56297 546821 56515
rect 546763 56233 546821 56239
rect 548391 56253 548449 56569
rect 549839 56260 549875 56498
rect 545129 56139 545135 56197
rect 545193 56139 545199 56197
rect 549831 56254 549883 56260
rect 549831 56196 549883 56202
rect 548391 56189 548449 56195
<< via1 >>
rect 265195 656552 265674 657031
rect 246223 653625 247829 655231
rect 321112 656552 321591 657031
rect 338957 653625 340563 655231
rect 560291 609925 560669 610303
rect 561263 609913 561641 610291
rect 72802 597575 72870 597643
rect 72744 595947 72812 596015
rect 76475 593643 76596 593764
rect 265195 566552 265674 567031
rect 246223 563625 247829 565231
rect 321112 566552 321591 567031
rect 338957 563625 340563 565231
rect 532586 522710 532670 522794
rect 532510 520206 532594 520290
rect 530211 501603 530297 501689
rect 530697 501161 530783 501247
rect 544533 488174 544619 488260
rect 542134 481542 542186 481594
rect 541952 480616 542004 480668
rect 265195 476552 265674 477031
rect 246223 473625 247829 475231
rect 321112 476552 321591 477031
rect 338957 473625 340563 475231
rect 52785 426798 52859 426872
rect 52877 426508 52951 426582
rect 52894 426023 53094 426223
rect 53035 425596 53109 425670
rect 53043 425314 53117 425388
rect 53035 425042 53109 425116
rect 53034 424701 53234 424901
rect 53034 424396 53234 424596
rect 34446 423301 34646 423501
rect 33750 423001 33950 423201
rect 33034 422701 33234 422901
rect 32362 422401 32562 422601
rect 37908 422101 38108 422301
rect 467308 388495 467444 388631
rect 467298 387792 467434 387928
rect 265195 386552 265674 387031
rect 246223 383625 247829 385231
rect 321112 386552 321591 387031
rect 467912 386128 468048 386264
rect 338957 383625 340563 385231
rect 468168 385111 468304 385247
rect 478342 383195 478416 383269
rect 461118 382157 461170 382209
rect 458196 381134 458332 381270
rect 486382 380907 486434 380959
rect 477002 379174 477054 379226
rect 488527 378502 488621 378596
rect 483683 378274 483777 378368
rect 487669 377992 487763 378086
rect 459335 377587 459589 377841
rect 459531 377189 459821 377479
rect 501381 376821 501711 377151
rect 459784 376009 460196 376421
rect 500454 375466 500534 375546
rect 502392 375466 502472 375546
rect 518984 375466 519064 375546
rect 459865 374677 460299 375111
rect 553602 373108 556478 376077
rect 556478 373108 556571 376077
rect 520746 372854 520826 372934
rect 442634 371062 443287 371715
rect 441444 367479 442145 368180
rect 520840 367864 520920 367944
rect 439833 364753 439963 364883
rect 577998 360764 580967 363733
rect 439337 347585 439555 347803
rect 483026 349242 483162 349378
rect 483044 348922 483180 349058
rect 483044 348584 483180 348720
rect 483078 348230 483214 348366
rect 483094 347960 483230 348096
rect 483128 347706 483264 347842
rect 483178 347436 483314 347572
rect 483212 347166 483348 347302
rect 38117 340170 38169 340222
rect 438563 329928 438742 330107
rect 519754 313890 519834 313970
rect 519594 313436 519674 313516
rect 519434 313084 519514 313164
rect 519274 312696 519354 312776
rect 519054 312150 519134 312230
rect 518894 311580 518974 311660
rect 518734 311150 518814 311230
rect 518574 310612 518654 310692
rect 265195 296552 265674 297031
rect 246223 293625 247829 295231
rect 321112 296552 321591 297031
rect 338957 293625 340563 295231
rect 265195 206552 265674 207031
rect 246223 203625 247829 205231
rect 321112 206552 321591 207031
rect 338957 203625 340563 205231
rect 552198 170290 552369 170461
rect 535443 152667 535501 152725
rect 537071 152435 537129 152493
rect 538699 152285 538757 152343
rect 540327 152121 540385 152179
rect 541955 151967 542013 152025
rect 543583 151729 543641 151787
rect 545211 151575 545269 151633
rect 546839 151417 546897 151475
rect 43657 131168 44035 131546
rect 43661 128787 44039 129165
rect 265195 116552 265674 117031
rect 246223 113625 247829 115231
rect 321112 116552 321591 117031
rect 338957 113625 340563 115231
rect 40028 58154 40164 59508
rect 536995 56451 537053 56509
rect 538623 56327 538681 56385
rect 540251 56349 540309 56407
rect 541879 56331 541937 56389
rect 543507 56267 543565 56325
rect 546763 56239 546821 56297
rect 545135 56139 545193 56197
rect 548391 56195 548449 56253
rect 549831 56202 549883 56254
<< metal2 >>
rect 137446 656216 138173 657462
rect 139419 657031 266022 657462
rect 139419 656552 265195 657031
rect 265674 656552 266022 657031
rect 139419 656216 266022 656552
rect 320764 657031 445405 657462
rect 320764 656552 321112 657031
rect 321591 656552 445405 657031
rect 320764 656216 445405 656552
rect 446651 656216 447266 657462
rect 246217 655062 246223 655231
rect 129998 653816 130007 655062
rect 131253 653816 246223 655062
rect 246217 653625 246223 653816
rect 247829 655062 247835 655231
rect 338951 655062 338957 655231
rect 247829 653816 248072 655062
rect 338714 653816 338957 655062
rect 247829 653625 247835 653816
rect 338951 653625 338957 653816
rect 340563 655062 340569 655231
rect 340563 653816 453593 655062
rect 454839 653816 454848 655062
rect 340563 653625 340569 653816
rect 279035 643726 282767 643786
rect 72802 597643 72870 597649
rect 72870 597575 76184 597643
rect 72802 597569 72870 597575
rect 72744 596015 72812 596021
rect 72812 595947 76024 596015
rect 72744 595941 72812 595947
rect 69966 563706 70006 566176
rect 70090 563830 70130 566176
rect 70206 563946 70246 566176
rect 70326 564066 70366 566176
rect 72558 564810 72598 566182
rect 72678 564930 72718 566182
rect 72798 565050 72838 566182
rect 72918 565170 72958 566182
rect 72918 565130 75864 565170
rect 72798 565010 75704 565050
rect 72678 564890 75484 564930
rect 72558 564770 75324 564810
rect 70326 564065 75110 564066
rect 70326 564026 75164 564065
rect 70206 563945 74944 563946
rect 70206 563906 75004 563945
rect 70090 563829 74746 563830
rect 70090 563790 74784 563829
rect 69966 563705 74554 563706
rect 69966 563666 74624 563705
rect 12150 509342 12220 510596
rect 12290 509502 12360 510596
rect 12430 509662 12500 510596
rect 12570 509822 12640 510596
rect 12570 509752 22284 509822
rect 12430 509592 22124 509662
rect 12290 509432 21964 509502
rect 12150 509272 21804 509342
rect 12150 466142 12220 467396
rect 12290 466302 12360 467396
rect 12430 466462 12500 467396
rect 12570 466622 12640 467396
rect 12570 466552 21284 466622
rect 12430 466392 21124 466462
rect 12290 466232 20964 466302
rect 12150 466072 20804 466142
rect 12150 422942 12220 424196
rect 12290 423102 12360 424196
rect 12430 423262 12500 424196
rect 12570 423422 12640 424196
rect 12570 423352 20284 423422
rect 12430 423192 20124 423262
rect 12290 423032 19964 423102
rect 12150 422872 19804 422942
rect 12150 379742 12220 380996
rect 12290 379902 12360 380996
rect 12430 380062 12500 380996
rect 12570 380222 12640 380996
rect 12570 380152 19284 380222
rect 12430 379992 19124 380062
rect 12290 379832 18964 379902
rect 12150 379672 18804 379742
rect 12150 336542 12220 337796
rect 12290 336702 12360 337796
rect 12430 336862 12500 337796
rect 12570 337022 12640 337796
rect 12570 336952 18284 337022
rect 12430 336792 18124 336862
rect 12290 336632 17964 336702
rect 12150 336472 17804 336542
rect 12150 293342 12220 294596
rect 12290 293502 12360 294596
rect 12430 293662 12500 294596
rect 12570 293822 12640 294596
rect 12570 293752 17284 293822
rect 12430 293592 17124 293662
rect 12290 293432 16964 293502
rect 12150 293272 16804 293342
rect 12150 250142 12220 251396
rect 12290 250302 12360 251396
rect 12430 250462 12500 251396
rect 12570 250622 12640 251396
rect 12570 250552 16284 250622
rect 12430 250392 16124 250462
rect 12290 250232 15964 250302
rect 12150 250072 15804 250142
rect 12714 120542 12784 123814
rect 12854 120702 12924 123814
rect 12994 120862 13064 123814
rect 13134 121022 13204 123814
rect 13134 120952 15284 121022
rect 12994 120792 15124 120862
rect 12854 120632 14964 120702
rect 12714 120472 14804 120542
rect 12714 77342 12784 80558
rect 12854 77502 12924 80558
rect 12994 77662 13064 80558
rect 13134 77822 13204 80558
rect 13134 77752 14284 77822
rect 12994 77592 14124 77662
rect 12854 77432 13964 77502
rect 12714 77272 13804 77342
rect 12714 2079 12784 37490
rect 12714 1964 12784 2009
rect 12854 2247 12924 37490
rect 12854 1964 12924 2177
rect 12994 2407 13064 37490
rect 12994 1964 13064 2337
rect 13134 2563 13204 37490
rect 13734 2723 13804 77272
rect 13734 2618 13804 2653
rect 13894 2883 13964 77432
rect 13894 2618 13964 2813
rect 14054 3043 14124 77592
rect 14054 2618 14124 2973
rect 14214 3199 14284 77752
rect 14734 3363 14804 120472
rect 14734 3244 14804 3293
rect 14894 3519 14964 120632
rect 14894 3244 14964 3449
rect 15054 3685 15124 120792
rect 15054 3244 15124 3615
rect 15214 3841 15284 120952
rect 15734 3999 15804 250072
rect 15734 3870 15804 3929
rect 15894 4167 15964 250232
rect 15894 3870 15964 4097
rect 16054 4327 16124 250392
rect 16054 3870 16124 4257
rect 16214 4489 16284 250552
rect 16734 4637 16804 293272
rect 16734 4536 16804 4567
rect 16894 4799 16964 293432
rect 16894 4536 16964 4729
rect 17054 4963 17124 293592
rect 17054 4536 17124 4893
rect 17214 5123 17284 293752
rect 17734 5281 17804 336472
rect 17734 5172 17804 5211
rect 17894 5443 17964 336632
rect 17894 5172 17964 5373
rect 18054 5607 18124 336792
rect 18054 5172 18124 5537
rect 18214 5763 18284 336952
rect 18734 5919 18804 379672
rect 18734 5798 18804 5849
rect 18894 6083 18964 379832
rect 18894 5798 18964 6013
rect 19054 6247 19124 379992
rect 19054 5798 19124 6177
rect 19214 6403 19284 380152
rect 19734 6563 19804 422872
rect 19734 6462 19804 6493
rect 19894 6725 19964 423032
rect 19894 6462 19964 6655
rect 20054 6885 20124 423192
rect 20054 6462 20124 6815
rect 20214 7045 20284 423352
rect 20734 7203 20804 466072
rect 20734 7080 20804 7133
rect 20894 7361 20964 466232
rect 20894 7080 20964 7291
rect 21054 7521 21124 466392
rect 21054 7080 21124 7451
rect 21214 7683 21284 466552
rect 21734 7845 21804 509272
rect 21734 7734 21804 7775
rect 21894 8005 21964 509432
rect 21894 7734 21964 7935
rect 22054 8167 22124 509592
rect 22054 7734 22124 8097
rect 22214 8323 22284 509752
rect 28406 496773 33694 497410
rect 28406 437437 29043 496773
rect 32420 496260 32488 496269
rect 32488 496192 33610 496260
rect 51168 496202 70696 496286
rect 70780 496202 70789 496286
rect 32420 496183 32488 496192
rect 30857 494838 30866 495378
rect 31406 494838 34087 495378
rect 32705 494100 32714 494160
rect 32774 494100 33610 494160
rect 31026 493286 31594 493298
rect 31026 492746 31040 493286
rect 31580 492746 34080 493286
rect 31026 492736 31594 492746
rect 32714 491644 74464 491646
rect 32707 491588 32716 491644
rect 32772 491588 74464 491644
rect 32714 491586 74464 491588
rect 32425 491500 32483 491504
rect 32420 491495 74304 491500
rect 32420 491437 32425 491495
rect 32483 491437 74304 491495
rect 32420 491432 74304 491437
rect 32425 491428 32483 491432
rect 34415 468680 34669 468684
rect 34410 468675 34674 468680
rect 34410 468421 34415 468675
rect 34669 468421 34674 468675
rect 33711 467974 33965 467978
rect 28406 437183 28647 437437
rect 28901 437183 29043 437437
rect 28406 436928 29043 437183
rect 33706 467969 33970 467974
rect 33706 467715 33711 467969
rect 33965 467715 33970 467969
rect 32303 424774 32557 424778
rect 32298 424769 32562 424774
rect 32298 424515 32303 424769
rect 32557 424515 32562 424769
rect 32298 422601 32562 424515
rect 33706 423201 33970 467715
rect 34410 423501 34674 468421
rect 52785 426872 52859 426878
rect 52859 426798 74084 426872
rect 52785 426792 52859 426798
rect 52877 426582 52951 426588
rect 52951 426508 73924 426582
rect 52877 426502 52951 426508
rect 52894 426223 53094 426229
rect 53094 426023 55450 426223
rect 55650 426023 55659 426223
rect 52894 426017 53094 426023
rect 53035 425670 53109 425676
rect 53109 425596 73764 425670
rect 53035 425590 53109 425596
rect 53043 425388 53117 425394
rect 53117 425314 73604 425388
rect 53043 425308 53117 425314
rect 53035 425116 53109 425122
rect 73314 425116 73384 425118
rect 53109 425042 73384 425116
rect 53035 425036 53109 425042
rect 53034 424901 53234 424907
rect 53234 424701 55426 424901
rect 55626 424701 55635 424901
rect 53034 424695 53234 424701
rect 53034 424596 53234 424602
rect 53234 424396 55428 424596
rect 55628 424396 55637 424596
rect 53034 424390 53234 424396
rect 34410 423301 34446 423501
rect 34646 423301 34674 423501
rect 34410 423246 34674 423301
rect 33706 423001 33750 423201
rect 33950 423001 33970 423201
rect 32962 422901 33226 422988
rect 33706 422940 33970 423001
rect 32962 422701 33034 422901
rect 33234 422701 33240 422901
rect 32298 422401 32362 422601
rect 32562 422401 32568 422601
rect 32298 422316 32562 422401
rect 32962 381569 33226 422701
rect 37908 422301 38108 422307
rect 37908 412914 38108 422101
rect 37908 412705 38108 412714
rect 32962 381315 32967 381569
rect 33221 381315 33226 381569
rect 32962 381310 33226 381315
rect 32967 381306 33221 381310
rect 23112 350808 23212 350817
rect 23112 332132 23212 350708
rect 38111 340170 38117 340222
rect 38169 340170 73224 340222
rect 36526 334472 40087 334978
rect 40593 334472 40602 334978
rect 36895 333578 40079 334060
rect 40561 333578 40570 334060
rect 23112 332032 25136 332132
rect 38766 331999 38866 332008
rect 36448 331899 38766 331999
rect 23112 331797 25136 331897
rect 38766 331890 38866 331899
rect 23124 307520 23224 331797
rect 24323 331339 24332 331439
rect 24432 331339 25368 331439
rect 23115 307420 23124 307520
rect 23224 307420 23233 307520
rect 40653 285265 42243 285274
rect 40653 275680 42243 283675
rect 44103 277951 45693 277970
rect 44103 276361 45657 277951
rect 47247 276361 47256 277951
rect 44103 275680 45693 276361
rect 39313 224282 39975 224305
rect 39313 223396 40406 224282
rect 39312 223387 40406 223396
rect 39964 222735 40406 223387
rect 39312 222730 40406 222735
rect 39312 222726 39964 222730
rect 40938 219528 41008 224321
rect 41298 219688 41368 224321
rect 41658 219848 41728 224295
rect 42078 220068 42148 224311
rect 42438 220228 42508 224343
rect 42798 220388 42868 224311
rect 43158 220548 43228 224315
rect 43578 220768 43648 224315
rect 43938 220928 44008 224359
rect 44298 221088 44368 224295
rect 44658 221248 44728 224289
rect 45078 221468 45148 224305
rect 45458 221628 45528 224311
rect 46119 224204 47252 224310
rect 46106 223542 61931 224204
rect 62593 223542 62602 224204
rect 45938 222730 45947 223392
rect 46609 222730 61877 223392
rect 62539 222730 62548 223392
rect 45458 221558 73064 221628
rect 45078 221398 72904 221468
rect 44658 221178 72684 221248
rect 44298 221018 72524 221088
rect 43938 220858 72364 220928
rect 43578 220698 72204 220768
rect 43158 220478 71984 220548
rect 42798 220318 71824 220388
rect 42438 220158 71664 220228
rect 42078 219998 71504 220068
rect 41658 219778 71284 219848
rect 41298 219618 71124 219688
rect 40938 219458 70964 219528
rect 41602 132506 44023 133617
rect 45134 132506 45143 133617
rect 43657 131546 44035 131552
rect 44035 131168 50123 131546
rect 50501 131168 50510 131546
rect 43657 131162 44035 131168
rect 42543 130806 42645 130810
rect 41848 130801 42650 130806
rect 41848 130699 42543 130801
rect 42645 130699 42650 130801
rect 41848 130694 42650 130699
rect 42543 130690 42645 130694
rect 41846 129804 70804 129872
rect 43661 129165 44039 129171
rect 44039 128787 50097 129165
rect 50475 128787 50484 129165
rect 43661 128781 44039 128787
rect 41480 126745 44572 127856
rect 45683 126745 45692 127856
rect 41188 59528 42568 59532
rect 40010 59523 42573 59528
rect 40010 59508 41188 59523
rect 40010 58154 40028 59508
rect 40164 58154 41188 59508
rect 40010 58143 41188 58154
rect 42568 58143 42573 59523
rect 40010 58138 42573 58143
rect 41188 58134 42568 58138
rect 42439 57258 42509 57267
rect 42424 57188 42439 57250
rect 42509 57188 42536 57250
rect 42424 9543 42536 57188
rect 42424 9441 42429 9543
rect 42531 9441 42536 9543
rect 42424 9436 42536 9441
rect 42732 57078 42844 57094
rect 42732 57008 42745 57078
rect 42815 57008 42844 57078
rect 42429 9432 42531 9436
rect 42732 9156 42844 57008
rect 42732 9147 42845 9156
rect 42732 9045 42743 9147
rect 42732 9036 42845 9045
rect 42732 9033 42844 9036
rect 70734 8483 70804 129804
rect 70734 8370 70804 8413
rect 70894 8643 70964 219458
rect 70894 8370 70964 8573
rect 71054 8803 71124 219618
rect 71054 8370 71124 8733
rect 71214 8963 71284 219778
rect 71434 9121 71504 219998
rect 71434 9014 71504 9051
rect 71594 9285 71664 220158
rect 71594 9014 71664 9215
rect 71754 9445 71824 220318
rect 71754 9014 71824 9375
rect 71914 9607 71984 220478
rect 72134 9765 72204 220698
rect 72134 9650 72204 9695
rect 72294 9925 72364 220858
rect 72294 9650 72364 9855
rect 72454 10085 72524 221018
rect 72454 9650 72524 10015
rect 72614 10243 72684 221178
rect 72834 10405 72904 221398
rect 72834 10286 72904 10335
rect 72994 10565 73064 221558
rect 72994 10286 73064 10495
rect 73154 10723 73224 340170
rect 73154 10286 73224 10653
rect 73314 10883 73384 425042
rect 73534 11047 73604 425314
rect 73534 10922 73604 10977
rect 73694 11201 73764 425596
rect 73694 10922 73764 11131
rect 73854 11363 73924 426508
rect 73854 10922 73924 11293
rect 74014 11523 74084 426798
rect 74234 11681 74304 491432
rect 74234 11576 74304 11611
rect 74394 11845 74464 491586
rect 74394 11576 74464 11775
rect 74554 12003 74624 563666
rect 74554 11576 74624 11933
rect 74714 12161 74784 563790
rect 74934 12325 75004 563906
rect 74934 12212 75004 12255
rect 75094 12481 75164 564026
rect 75094 12212 75164 12411
rect 75254 12643 75324 564770
rect 75254 12212 75324 12573
rect 75414 12803 75484 564890
rect 75634 12963 75704 565010
rect 75634 12838 75704 12893
rect 75794 13121 75864 565130
rect 75794 12838 75864 13051
rect 75954 13283 76024 595947
rect 75954 12838 76024 13213
rect 76114 13447 76184 597575
rect 76475 593764 76596 593770
rect 76596 593643 87042 593764
rect 76475 593637 76596 593643
rect 86921 591465 87042 593643
rect 86921 591344 126893 591465
rect 127014 591344 127023 591465
rect 137828 566216 138287 567462
rect 139533 567031 266022 567462
rect 139533 566552 265195 567031
rect 265674 566552 266022 567031
rect 139533 566216 266022 566552
rect 246217 565062 246223 565231
rect 129998 563816 130007 565062
rect 131253 563816 246223 565062
rect 246217 563625 246223 563816
rect 247829 565062 247835 565231
rect 247829 563816 248072 565062
rect 247829 563625 247835 563816
rect 279035 553726 282487 553786
rect 130489 520258 130498 520554
rect 130794 520258 130803 520554
rect 138454 519191 138463 519501
rect 138773 519191 138782 519501
rect 137676 476216 138401 477462
rect 139647 477031 266022 477462
rect 139647 476552 265195 477031
rect 265674 476552 266022 477031
rect 139647 476216 266022 476552
rect 246217 475062 246223 475231
rect 130150 473816 130159 475062
rect 131405 473816 246223 475062
rect 246217 473625 246223 473816
rect 247829 475062 247835 475231
rect 247829 473816 248072 475062
rect 247829 473625 247835 473816
rect 279035 463726 282207 463786
rect 137676 386216 138267 387462
rect 139513 387031 266022 387462
rect 139513 386552 265195 387031
rect 265674 386552 266022 387031
rect 139513 386216 266022 386552
rect 246217 385062 246223 385231
rect 130150 383816 130159 385062
rect 131405 383816 246223 385062
rect 246217 383625 246223 383816
rect 247829 385062 247835 385231
rect 247829 383816 248072 385062
rect 247829 383625 247835 383816
rect 279035 373726 281927 373786
rect 137446 296216 138115 297462
rect 139361 297031 266022 297462
rect 139361 296552 265195 297031
rect 265674 296552 266022 297031
rect 139361 296216 266022 296552
rect 246217 295062 246223 295231
rect 129920 293816 129929 295062
rect 131175 293816 246223 295062
rect 246217 293625 246223 293816
rect 247829 295062 247835 295231
rect 247829 293816 248072 295062
rect 247829 293625 247835 293816
rect 279035 283726 281647 283786
rect 137598 206216 138191 207462
rect 139437 207031 266022 207462
rect 139437 206552 265195 207031
rect 265674 206552 266022 207031
rect 139437 206216 266022 206552
rect 246217 205062 246223 205231
rect 130150 203816 130159 205062
rect 131405 203816 246223 205062
rect 246217 203625 246223 203816
rect 247829 205062 247835 205231
rect 247829 203816 248072 205062
rect 247829 203625 247835 203816
rect 279035 193726 281367 193786
rect 137446 116216 138173 117462
rect 139419 117031 266022 117462
rect 139419 116552 265195 117031
rect 265674 116552 266022 117031
rect 139419 116216 266022 116552
rect 246217 115062 246223 115231
rect 129998 113816 130007 115062
rect 131253 113816 246223 115062
rect 246217 113625 246223 113816
rect 247829 115062 247835 115231
rect 247829 113816 248072 115062
rect 247829 113625 247835 113816
rect 279035 103726 281087 103786
rect 76114 12838 76184 13377
rect 253067 13445 253198 13469
rect 253067 13374 253096 13445
rect 253167 13374 253198 13445
rect 251883 13285 252014 13311
rect 251883 13214 251904 13285
rect 251975 13214 252014 13285
rect 249533 13125 249655 13145
rect 249533 13054 249554 13125
rect 249625 13054 249655 13125
rect 248349 12965 248471 12981
rect 248349 12894 248370 12965
rect 248441 12894 248471 12965
rect 75414 12212 75484 12733
rect 246011 12811 246101 12820
rect 244827 12651 244917 12660
rect 242475 12497 242565 12506
rect 241291 12335 241381 12344
rect 74714 11576 74784 12091
rect 238927 12173 239017 12182
rect 237743 12011 237833 12020
rect 235362 11854 235462 11863
rect 234178 11696 234278 11708
rect 74014 10922 74084 11453
rect 231814 11542 231914 11551
rect 230630 11384 230730 11393
rect 228288 11224 228388 11233
rect 227104 11060 227204 11069
rect 73314 10286 73384 10813
rect 224740 10900 224840 10909
rect 223556 10742 223656 10751
rect 221202 10584 221302 10593
rect 220018 10422 220118 10431
rect 72614 9650 72684 10173
rect 217644 10245 217744 10276
rect 217644 10174 217658 10245
rect 217729 10174 217744 10245
rect 216476 10090 216547 10094
rect 216460 10085 216560 10090
rect 216460 10014 216476 10085
rect 216547 10014 216560 10085
rect 214129 9920 214198 9929
rect 212945 9758 213014 9767
rect 71914 9014 71984 9537
rect 210577 9596 210646 9605
rect 209393 9438 209462 9447
rect 207019 9292 207088 9301
rect 205835 9134 205904 9143
rect 71214 8370 71284 8893
rect 203478 8960 203538 8969
rect 203478 8891 203538 8900
rect 202294 8811 202353 8859
rect 202294 8802 202354 8811
rect 202294 8733 202354 8742
rect 199920 8661 200010 8670
rect 198736 8491 198826 8532
rect 22214 7734 22284 8253
rect 196359 8339 196449 8351
rect 195175 8173 195265 8182
rect 192827 7991 192897 8029
rect 191643 7849 191713 7868
rect 21214 7080 21284 7613
rect 189287 7694 189368 7716
rect 188103 7520 188184 7554
rect 185747 7372 185828 7392
rect 184563 7218 184644 7238
rect 20214 6462 20284 6975
rect 182183 7050 182264 7080
rect 180999 6896 181080 6912
rect 178632 6732 178713 6762
rect 177448 6574 177529 6596
rect 19214 5798 19284 6333
rect 175093 6408 175174 6438
rect 173909 6248 173990 6272
rect 171566 6094 171647 6130
rect 170382 5930 170463 5958
rect 18214 5172 18284 5693
rect 168002 5768 168083 5798
rect 166818 5608 166899 5636
rect 164457 5446 164538 5468
rect 163273 5302 163354 5320
rect 17214 4536 17284 5053
rect 160918 5124 160999 5150
rect 159734 4956 159815 4990
rect 157360 4806 157441 4838
rect 156176 4652 156257 4692
rect 16214 3870 16284 4419
rect 153808 4488 153889 4512
rect 152624 4334 152705 4356
rect 150282 4170 150363 4184
rect 149098 4008 149179 4032
rect 15214 3244 15284 3771
rect 146724 3852 146805 3866
rect 145540 3694 145621 3716
rect 143191 3534 143272 3554
rect 142007 3368 142088 3404
rect 14214 2618 14284 3129
rect 139633 3216 139714 3238
rect 138449 3050 138530 3080
rect 136088 2900 136169 2938
rect 134904 2728 134985 2756
rect 13134 1964 13204 2493
rect 132555 2562 132636 2598
rect 131371 2406 131452 2432
rect 129002 2260 129083 2274
rect 127818 2088 127899 2104
rect 1324 800 1436 1280
rect 2506 800 2618 1280
rect 3688 800 3800 1280
rect 4870 800 4982 1280
rect 6052 800 6164 1280
rect 7234 800 7346 1280
rect 8416 800 8528 1280
rect 9598 800 9710 1280
rect 10780 800 10892 1280
rect 11962 800 12074 1280
rect 13144 800 13256 1280
rect 14326 800 14438 1280
rect 15508 800 15620 1280
rect 16690 800 16802 1280
rect 17872 800 17984 1280
rect 19054 800 19166 1280
rect 20236 800 20348 1280
rect 21418 800 21530 1280
rect 22600 800 22712 1280
rect 23782 800 23894 1280
rect 24964 800 25076 1280
rect 26146 800 26258 1280
rect 27328 800 27440 1280
rect 28510 800 28622 1280
rect 29692 800 29804 1280
rect 30874 800 30986 1280
rect 32056 800 32168 1280
rect 33238 800 33350 1280
rect 34420 800 34532 1280
rect 35602 800 35714 1280
rect 36784 800 36896 1280
rect 37966 800 38078 1280
rect 39148 800 39260 1280
rect 40330 800 40442 1280
rect 41512 800 41624 1280
rect 42694 800 42806 1280
rect 43876 800 43988 1280
rect 45058 800 45170 1280
rect 46240 800 46352 1280
rect 47422 800 47534 1280
rect 48604 800 48716 1280
rect 49786 800 49898 1280
rect 50968 800 51080 1280
rect 52150 800 52262 1280
rect 53332 800 53444 1280
rect 54514 800 54626 1280
rect 55696 800 55808 1280
rect 56878 800 56990 1280
rect 58060 800 58172 1280
rect 59242 800 59354 1280
rect 60424 800 60536 1280
rect 61606 800 61718 1280
rect 62788 800 62900 1280
rect 63970 800 64082 1280
rect 65152 800 65264 1280
rect 66334 800 66446 1280
rect 67516 800 67628 1280
rect 68698 800 68810 1280
rect 69880 800 69992 1280
rect 71062 800 71174 1280
rect 72244 800 72356 1280
rect 73426 800 73538 1280
rect 74608 800 74720 1280
rect 75790 800 75902 1280
rect 76972 800 77084 1280
rect 78154 800 78266 1280
rect 79336 800 79448 1280
rect 80518 800 80630 1280
rect 81700 800 81812 1280
rect 82882 800 82994 1280
rect 84064 800 84176 1280
rect 85246 800 85358 1280
rect 86428 800 86540 1280
rect 87610 800 87722 1280
rect 88792 800 88904 1280
rect 89974 800 90086 1280
rect 91156 800 91268 1280
rect 92338 800 92450 1280
rect 93520 800 93632 1280
rect 94702 800 94814 1280
rect 95884 800 95996 1280
rect 97066 800 97178 1280
rect 98248 800 98360 1280
rect 99430 800 99542 1280
rect 100612 800 100724 1280
rect 101794 800 101906 1280
rect 102976 800 103088 1280
rect 104158 800 104270 1280
rect 105340 800 105452 1280
rect 106522 800 106634 1280
rect 107704 800 107816 1280
rect 108886 800 108998 1280
rect 110068 800 110180 1279
rect 111250 800 111362 1280
rect 112432 800 112544 1280
rect 113614 800 113726 1280
rect 114796 800 114908 1280
rect 115978 800 116090 1280
rect 117160 800 117272 1280
rect 118342 800 118454 1280
rect 119524 800 119636 1280
rect 120706 800 120818 1280
rect 121888 800 122000 1280
rect 123070 800 123182 1280
rect 124252 800 124364 1280
rect 125434 800 125546 1280
rect 126616 800 126728 1280
rect 127818 1258 127899 2007
rect 129002 1280 129083 2179
rect 131371 1280 131452 2325
rect 132555 1280 132636 2481
rect 134904 1280 134985 2647
rect 136088 1280 136169 2819
rect 138449 1280 138530 2969
rect 127798 800 127910 1258
rect 128980 800 129092 1280
rect 130162 800 130274 1280
rect 129002 0 129083 800
rect 131344 0 131456 1280
rect 132526 800 132638 1280
rect 133708 800 133820 1280
rect 132555 0 132636 800
rect 134890 0 135002 1280
rect 136072 800 136184 1280
rect 137254 800 137366 1280
rect 136088 0 136169 800
rect 138436 0 138548 1280
rect 139633 1279 139714 3135
rect 142007 1280 142088 3287
rect 139618 800 139730 1279
rect 140800 800 140912 1279
rect 139633 0 139714 800
rect 141982 0 142094 1280
rect 143191 1279 143272 3453
rect 145540 1280 145621 3613
rect 145528 1279 145640 1280
rect 146724 1279 146805 3771
rect 149098 1280 149179 3927
rect 143164 800 143276 1279
rect 144346 800 144458 1279
rect 145528 1178 145648 1279
rect 143191 0 143272 800
rect 145528 0 145640 1178
rect 146710 800 146822 1279
rect 147892 800 148004 1279
rect 146724 0 146805 800
rect 149074 0 149186 1280
rect 150282 1279 150363 4089
rect 152624 1280 152705 4253
rect 150256 800 150368 1279
rect 151438 800 151550 1279
rect 152614 1096 152732 1280
rect 153808 1279 153889 4407
rect 156176 1280 156257 4571
rect 150282 0 150363 800
rect 152620 0 152732 1096
rect 153802 800 153914 1279
rect 154984 800 155096 1279
rect 153808 0 153889 800
rect 156166 0 156278 1280
rect 157360 1279 157441 4725
rect 159734 1280 159815 4875
rect 159712 1279 159824 1280
rect 160918 1279 160999 5043
rect 163273 1280 163354 5221
rect 163258 1279 163370 1280
rect 164457 1279 164538 5365
rect 166818 1280 166899 5527
rect 166804 1279 166916 1280
rect 168002 1279 168083 5687
rect 170382 1280 170463 5849
rect 170350 1279 170464 1280
rect 171566 1279 171647 6013
rect 173909 1280 173990 6167
rect 157348 800 157460 1279
rect 158530 800 158642 1279
rect 159712 1152 159836 1279
rect 157360 0 157441 800
rect 159712 0 159824 1152
rect 160894 800 161006 1279
rect 162076 800 162188 1279
rect 163258 1108 163374 1279
rect 160918 0 160999 800
rect 163258 0 163370 1108
rect 164440 800 164552 1279
rect 165622 800 165734 1279
rect 166804 1140 166922 1279
rect 164457 0 164538 800
rect 166804 0 166916 1140
rect 167986 800 168098 1279
rect 169168 800 169280 1279
rect 170348 1130 170464 1279
rect 170350 1112 170464 1130
rect 171532 1112 171647 1279
rect 168002 0 168083 800
rect 170350 0 170462 1112
rect 171532 800 171644 1112
rect 172714 800 172826 1279
rect 173896 0 174008 1280
rect 175093 1279 175174 6327
rect 177448 1280 177529 6493
rect 175078 800 175190 1279
rect 176260 800 176372 1279
rect 175093 0 175174 800
rect 177442 0 177554 1280
rect 178632 1279 178713 6651
rect 180999 1280 181080 6815
rect 178624 800 178736 1279
rect 179806 800 179918 1279
rect 178632 0 178713 800
rect 180988 0 181100 1280
rect 182183 1279 182264 6969
rect 184563 1280 184644 7137
rect 182170 800 182282 1279
rect 183352 800 183464 1279
rect 182183 0 182264 800
rect 184534 0 184646 1280
rect 185747 1279 185828 7291
rect 188103 1280 188184 7439
rect 186929 1279 186987 1280
rect 185716 800 185828 1279
rect 186898 800 187010 1279
rect 185747 0 185828 800
rect 188080 0 188192 1280
rect 189287 1279 189368 7613
rect 191643 1280 191713 7779
rect 190445 1279 190547 1280
rect 189262 800 189374 1279
rect 190444 800 190556 1279
rect 191621 1141 191738 1280
rect 192827 1279 192897 7921
rect 195175 1280 195265 8083
rect 189287 0 189368 800
rect 191626 0 191738 1141
rect 192808 800 192920 1279
rect 193990 800 194102 1279
rect 192827 0 192897 800
rect 195172 0 195284 1280
rect 196359 1279 196449 8249
rect 198736 1280 198826 8401
rect 199920 1280 200010 8571
rect 202294 1280 202353 8733
rect 203478 1280 203537 8891
rect 205835 1280 205904 9065
rect 207019 1280 207088 9223
rect 209393 1280 209462 9369
rect 210577 1280 210646 9527
rect 212945 1280 213014 9689
rect 214129 1280 214198 9851
rect 216460 1280 216560 10014
rect 217644 1280 217744 10174
rect 220018 1280 220118 10322
rect 221202 1280 221302 10484
rect 223556 1280 223656 10642
rect 224740 1280 224840 10800
rect 227104 1280 227204 10960
rect 228288 1280 228388 11124
rect 230630 1280 230730 11284
rect 231814 1280 231914 11442
rect 234178 1280 234278 11596
rect 235362 1280 235462 11754
rect 237743 1280 237833 11921
rect 238927 1280 239017 12083
rect 241291 1280 241381 12245
rect 242475 1280 242565 12407
rect 244827 1280 244917 12561
rect 246011 1280 246101 12721
rect 248349 1280 248471 12894
rect 249533 1280 249655 13054
rect 251883 1280 252014 13214
rect 253067 1280 253198 13374
rect 280296 9936 280356 9945
rect 276749 9760 276809 9769
rect 273201 9610 273261 9619
rect 255461 1280 255583 1416
rect 256645 1280 256767 1416
rect 259000 1280 259100 1416
rect 260184 1280 260284 1416
rect 262570 1280 262630 1416
rect 263754 1280 263814 1416
rect 266118 1280 266178 1416
rect 269654 1280 269714 1508
rect 273201 1280 273261 9550
rect 276749 1280 276809 9700
rect 280296 1280 280356 9876
rect 281027 9588 281087 103726
rect 281307 9750 281367 193726
rect 281587 9912 281647 283726
rect 281867 10066 281927 373726
rect 282147 10228 282207 463726
rect 282427 10406 282487 553726
rect 282707 10544 282767 643726
rect 303962 643726 307687 643786
rect 282707 10475 282767 10484
rect 294486 10568 294546 10577
rect 282427 10337 282487 10346
rect 290938 10410 290998 10419
rect 282147 10159 282207 10168
rect 287391 10252 287451 10261
rect 281867 9997 281927 10006
rect 283843 10102 283903 10111
rect 281587 9843 281647 9852
rect 281307 9681 281367 9690
rect 281027 9519 281087 9528
rect 283843 1280 283903 10042
rect 287391 1280 287451 10192
rect 290938 1280 290998 10350
rect 294486 1280 294546 10508
rect 298033 9440 298093 9449
rect 298033 1280 298093 9380
rect 303962 9442 304022 643726
rect 538242 613613 538251 615607
rect 540245 613613 546564 615607
rect 558734 611592 583269 611666
rect 583343 611592 583352 611666
rect 558744 610762 559378 610836
rect 540996 606980 541059 608974
rect 543053 606980 546582 608974
rect 518034 605409 518114 605410
rect 559299 605409 559373 610762
rect 518034 605335 559373 605409
rect 560291 610303 560669 610309
rect 454025 592807 454034 593103
rect 454330 592807 454339 593103
rect 320764 567031 445481 567462
rect 320764 566552 321112 567031
rect 321591 566552 445481 567031
rect 320764 566216 445481 566552
rect 446727 566216 447342 567462
rect 338951 565062 338957 565231
rect 338714 563816 338957 565062
rect 338951 563625 338957 563816
rect 340563 565062 340569 565231
rect 340563 563816 453515 565062
rect 454761 563816 454770 565062
rect 340563 563625 340569 563816
rect 303962 9373 304022 9382
rect 304242 553726 307687 553786
rect 301569 9282 301629 9291
rect 301569 1280 301629 9222
rect 304242 9272 304302 553726
rect 445832 494877 445841 495187
rect 446151 494877 446160 495187
rect 454071 483040 454080 483336
rect 454376 483040 454385 483336
rect 320764 477031 445367 477462
rect 320764 476552 321112 477031
rect 321591 476552 445367 477031
rect 320764 476216 445367 476552
rect 446613 476216 447266 477462
rect 338951 475062 338957 475231
rect 338714 473816 338957 475062
rect 338951 473625 338957 473816
rect 340563 475062 340569 475231
rect 340563 473816 453439 475062
rect 454685 473816 454694 475062
rect 340563 473625 340569 473816
rect 304242 9203 304302 9212
rect 304522 463726 307687 463786
rect 304522 9118 304582 463726
rect 467308 388631 467444 388637
rect 467444 388495 517544 388631
rect 517680 388495 517689 388631
rect 467308 388489 467444 388495
rect 467298 387928 467434 387934
rect 467434 387792 517556 387928
rect 517692 387792 517701 387928
rect 467298 387786 467434 387792
rect 320764 387031 445481 387462
rect 320764 386552 321112 387031
rect 321591 386552 445481 387031
rect 320764 386216 445481 386552
rect 446727 386216 447342 387462
rect 467912 386264 468048 386270
rect 468048 386128 517688 386264
rect 517824 386128 517833 386264
rect 467912 386122 468048 386128
rect 468168 385247 468304 385253
rect 338951 385062 338957 385231
rect 338714 383816 338957 385062
rect 338951 383625 338957 383816
rect 340563 385062 340569 385231
rect 468304 385111 517526 385247
rect 517662 385111 517671 385247
rect 468168 385105 468304 385111
rect 340563 383816 453515 385062
rect 454761 383816 454770 385062
rect 340563 383625 340569 383816
rect 478336 383195 478342 383269
rect 478416 383195 516805 383269
rect 516879 383195 516888 383269
rect 451707 382200 451716 382213
rect 451702 382166 451716 382200
rect 451707 382153 451716 382166
rect 451776 382200 451785 382213
rect 461112 382200 461118 382209
rect 451776 382166 461118 382200
rect 451776 382153 451785 382166
rect 461112 382157 461118 382166
rect 461170 382157 461176 382209
rect 441444 381752 442145 381761
rect 439337 381475 439555 381484
rect 438563 381377 438742 381386
rect 304522 9049 304582 9058
rect 304802 373726 307687 373786
rect 304802 8956 304862 373726
rect 438563 330107 438742 381198
rect 439337 347803 439555 381257
rect 439824 381255 439833 381385
rect 439963 381255 439972 381385
rect 439833 364883 439963 381255
rect 441444 368180 442145 381051
rect 442634 381672 443287 381681
rect 458196 381270 458332 381276
rect 451214 381134 451236 381270
rect 451372 381134 458196 381270
rect 458196 381128 458332 381134
rect 442634 371715 443287 381019
rect 486370 380959 486468 380966
rect 486370 380907 486382 380959
rect 486434 380958 486468 380959
rect 506913 380958 506922 380963
rect 486434 380908 506922 380958
rect 486434 380907 486468 380908
rect 486370 380902 486468 380907
rect 506913 380903 506922 380908
rect 506982 380903 506991 380963
rect 476996 379174 477002 379226
rect 477054 379174 477060 379226
rect 477002 378840 477054 379174
rect 516870 378844 516930 378853
rect 477002 378788 516870 378840
rect 516870 378775 516930 378784
rect 488527 378596 488621 378602
rect 488621 378502 516821 378596
rect 516915 378502 516924 378596
rect 488527 378496 488621 378502
rect 483683 378368 483777 378374
rect 483777 378274 516881 378368
rect 516975 378274 516984 378368
rect 483683 378268 483777 378274
rect 487669 378086 487763 378092
rect 487763 377992 516953 378086
rect 517047 377992 517056 378086
rect 487669 377986 487763 377992
rect 459335 377841 459589 377847
rect 459260 377587 459335 377841
rect 459589 377751 462022 377756
rect 459589 377649 461915 377751
rect 462017 377649 462026 377751
rect 459589 377644 462022 377649
rect 459335 377581 459589 377587
rect 459531 377479 459821 377485
rect 459260 377189 459531 377479
rect 459821 377385 461302 377390
rect 459821 377283 461195 377385
rect 461297 377283 461306 377385
rect 459821 377278 461302 377283
rect 459531 377183 459821 377189
rect 501375 376821 501381 377151
rect 501711 376821 505921 377151
rect 506251 376821 506260 377151
rect 459784 376421 460196 376427
rect 450382 376009 450424 376421
rect 450836 376009 459784 376421
rect 459784 376003 460196 376009
rect 502392 375546 502472 375552
rect 500448 375466 500454 375546
rect 500534 375466 502392 375546
rect 502392 375460 502472 375466
rect 449312 375111 449774 375122
rect 459865 375111 460299 375117
rect 449312 374677 449325 375111
rect 449759 374677 459865 375111
rect 449312 374668 449774 374677
rect 459865 374671 460299 374677
rect 442634 371056 443287 371062
rect 441444 367473 442145 367479
rect 439833 364747 439963 364753
rect 483026 349378 483162 349384
rect 483162 349242 490958 349378
rect 491094 349242 491103 349378
rect 483026 349236 483162 349242
rect 483038 348922 483044 349058
rect 483180 348922 490906 349058
rect 491042 348922 491051 349058
rect 483044 348720 483180 348726
rect 490890 348720 491026 348729
rect 483180 348584 490890 348720
rect 483044 348578 483180 348584
rect 490890 348575 491026 348584
rect 490958 348366 491094 348375
rect 483072 348230 483078 348366
rect 483214 348230 490958 348366
rect 490958 348221 491094 348230
rect 483094 348096 483230 348102
rect 483230 347960 490822 348096
rect 490958 347960 490967 348096
rect 483094 347954 483230 347960
rect 483128 347842 483264 347848
rect 490822 347842 490958 347851
rect 439331 347585 439337 347803
rect 439555 347585 439561 347803
rect 483264 347706 490822 347842
rect 483128 347700 483264 347706
rect 490822 347697 490958 347706
rect 483172 347436 483178 347572
rect 483314 347436 490890 347572
rect 491026 347436 491035 347572
rect 483206 347166 483212 347302
rect 483348 347166 490940 347302
rect 491076 347166 491085 347302
rect 438563 329922 438742 329928
rect 320764 297031 445367 297462
rect 320764 296552 321112 297031
rect 321591 296552 445367 297031
rect 320764 296216 445367 296552
rect 446613 296216 447188 297462
rect 338951 295062 338957 295231
rect 338714 293816 338957 295062
rect 338951 293625 338957 293816
rect 340563 295062 340569 295231
rect 453707 295062 454953 295071
rect 340563 293816 453707 295062
rect 454953 293816 454962 295052
rect 340563 293625 340569 293816
rect 453707 293807 454953 293816
rect 305082 283726 307687 283786
rect 304793 8896 304802 8956
rect 304862 8896 304871 8956
rect 305082 8778 305142 283726
rect 320764 207031 445597 207462
rect 320764 206552 321112 207031
rect 321591 206552 445597 207031
rect 320764 206216 445597 206552
rect 446843 206216 447188 207462
rect 338951 205062 338957 205231
rect 338714 203816 338957 205062
rect 338951 203625 338957 203816
rect 340563 205062 340569 205231
rect 340563 203816 453325 205062
rect 454571 203816 454580 205062
rect 340563 203625 340569 203816
rect 305082 8709 305142 8718
rect 305362 193726 307687 193786
rect 305362 8632 305422 193726
rect 320764 117031 445481 117462
rect 320764 116552 321112 117031
rect 321591 116552 445481 117031
rect 320764 116216 445481 116552
rect 446727 116216 447188 117462
rect 338951 115062 338957 115231
rect 338714 113816 338957 115062
rect 338951 113625 338957 113816
rect 340563 115062 340569 115231
rect 340563 113816 453593 115062
rect 454839 113816 454848 115062
rect 340563 113625 340569 113816
rect 305642 103726 307687 103786
rect 305353 8572 305362 8632
rect 305422 8572 305431 8632
rect 305362 8563 305418 8572
rect 305642 8486 305702 103726
rect 448122 14678 448239 14687
rect 305642 8417 305702 8426
rect 306122 9128 306182 9137
rect 306122 7852 306182 9068
rect 305122 7792 306182 7852
rect 308682 8962 308742 8971
rect 305122 1280 305182 7792
rect 308682 1280 308742 8902
rect 312210 8810 312270 8819
rect 312210 1280 312270 8750
rect 315770 8660 315830 8669
rect 315770 1280 315830 8600
rect 319309 8484 319369 8493
rect 319309 1280 319369 8424
rect 322858 1280 322918 1918
rect 326397 1280 326457 1918
rect 329936 1280 329996 2566
rect 333496 1280 333556 2566
rect 337045 1280 337105 2804
rect 340584 1280 340644 2804
rect 344133 1280 344193 2804
rect 347693 1280 347753 2804
rect 351221 1280 351281 2804
rect 354767 1280 354827 2804
rect 358322 1280 358382 2804
rect 361844 1280 361904 2804
rect 365396 1280 365456 2804
rect 368961 1280 369021 2804
rect 372480 1280 372540 2804
rect 376051 1280 376111 2804
rect 379597 1280 379657 2804
rect 383149 1280 383209 2804
rect 386688 1280 386748 2804
rect 390233 1280 390293 2804
rect 393785 1280 393845 2804
rect 397343 1280 397403 2804
rect 400869 1280 400929 2804
rect 404410 1280 404470 2804
rect 407958 1280 408018 2804
rect 411506 1280 411566 2804
rect 415054 1280 415114 2804
rect 418602 1280 418662 2804
rect 422150 1280 422210 2804
rect 425698 1280 425758 2804
rect 196354 800 196466 1279
rect 197536 800 197648 1279
rect 196359 0 196449 800
rect 198718 0 198830 1280
rect 199900 800 200012 1280
rect 201082 800 201194 1280
rect 199920 0 200010 800
rect 202264 0 202376 1280
rect 203446 800 203558 1280
rect 204628 800 204740 1280
rect 203478 0 203537 800
rect 205810 0 205922 1280
rect 206992 800 207104 1280
rect 208174 800 208286 1280
rect 207019 0 207088 800
rect 209356 0 209468 1280
rect 210538 800 210650 1280
rect 211720 800 211832 1280
rect 212902 800 213014 1280
rect 214084 800 214198 1280
rect 215266 800 215378 1280
rect 210577 0 210646 800
rect 212910 0 213014 800
rect 214129 0 214198 800
rect 216448 0 216560 1280
rect 217630 800 217744 1280
rect 218812 800 218924 1280
rect 219994 1279 220118 1280
rect 221176 1279 221302 1280
rect 217644 0 217744 800
rect 219994 0 220106 1279
rect 221176 800 221288 1279
rect 222358 800 222470 1280
rect 223540 1279 223656 1280
rect 224722 1279 224840 1280
rect 223540 0 223652 1279
rect 224722 800 224834 1279
rect 225904 800 226016 1280
rect 227086 1279 227204 1280
rect 228268 1279 228388 1280
rect 227086 0 227198 1279
rect 228268 800 228380 1279
rect 229450 800 229562 1280
rect 230630 1279 230744 1280
rect 230632 0 230744 1279
rect 231814 800 231926 1280
rect 232996 800 233108 1280
rect 234178 0 234290 1280
rect 235360 800 235472 1280
rect 236542 800 236654 1280
rect 235362 0 235462 800
rect 237724 0 237836 1280
rect 238906 800 239018 1280
rect 240088 800 240200 1280
rect 238927 0 239017 800
rect 241270 0 241382 1280
rect 242452 800 242565 1280
rect 243634 800 243746 1280
rect 242475 0 242565 800
rect 244816 0 244928 1280
rect 245998 800 246110 1280
rect 247180 800 247292 1280
rect 246011 0 246101 800
rect 248362 0 248474 1280
rect 249544 800 249656 1280
rect 250726 800 250838 1280
rect 251908 0 252020 1280
rect 253090 800 253202 1280
rect 254272 800 254384 1280
rect 255454 0 255566 1280
rect 256636 800 256748 1280
rect 257818 800 257930 1280
rect 259000 0 259112 1280
rect 260182 800 260294 1280
rect 261364 800 261476 1280
rect 260184 0 260284 800
rect 262546 0 262658 1280
rect 263728 800 263840 1280
rect 264910 800 265022 1280
rect 263754 0 263814 800
rect 266092 0 266204 1280
rect 267274 800 267386 1280
rect 268456 800 268568 1280
rect 269638 1175 269752 1280
rect 269638 0 269750 1175
rect 270820 800 270932 1280
rect 272002 800 272114 1280
rect 273184 0 273296 1280
rect 274366 800 274478 1280
rect 275548 800 275660 1280
rect 276730 0 276842 1280
rect 277912 800 278024 1280
rect 279094 800 279206 1280
rect 280276 0 280388 1280
rect 281458 800 281570 1280
rect 282640 800 282752 1280
rect 283822 0 283934 1280
rect 285004 800 285116 1280
rect 286186 800 286298 1280
rect 287368 0 287480 1280
rect 288550 800 288662 1280
rect 289732 800 289844 1280
rect 290914 0 291026 1280
rect 292096 800 292208 1280
rect 293278 800 293390 1280
rect 294460 0 294572 1280
rect 295642 800 295754 1280
rect 296824 800 296936 1280
rect 298006 0 298118 1280
rect 299188 800 299300 1280
rect 300370 800 300482 1280
rect 301552 0 301664 1280
rect 302734 800 302846 1280
rect 303916 800 304028 1280
rect 305098 0 305210 1280
rect 306280 800 306392 1280
rect 307462 800 307574 1280
rect 308644 0 308756 1280
rect 309826 800 309938 1280
rect 311008 800 311120 1280
rect 312190 0 312302 1280
rect 313372 800 313484 1280
rect 314554 800 314666 1280
rect 315736 0 315848 1280
rect 316918 800 317030 1280
rect 318100 800 318212 1280
rect 319282 0 319394 1280
rect 320464 800 320576 1280
rect 321646 800 321758 1280
rect 322828 0 322940 1280
rect 324010 800 324122 1280
rect 325192 800 325304 1280
rect 326374 0 326486 1280
rect 327556 800 327668 1280
rect 328738 800 328850 1280
rect 329920 0 330032 1280
rect 331102 800 331214 1280
rect 332284 800 332396 1280
rect 333466 0 333578 1280
rect 334648 800 334760 1280
rect 335830 800 335942 1280
rect 337012 0 337124 1280
rect 338194 800 338306 1280
rect 339376 800 339488 1280
rect 340558 0 340670 1280
rect 341740 800 341852 1280
rect 342922 800 343034 1280
rect 344104 0 344216 1280
rect 345286 800 345398 1280
rect 346468 800 346580 1280
rect 347650 0 347762 1280
rect 348832 800 348944 1280
rect 350014 800 350126 1280
rect 351196 0 351308 1280
rect 352378 800 352490 1280
rect 353560 800 353672 1280
rect 354742 0 354854 1280
rect 355924 800 356036 1280
rect 357106 800 357218 1280
rect 358288 0 358400 1280
rect 359470 800 359582 1280
rect 360652 800 360764 1280
rect 361834 0 361946 1280
rect 363016 800 363128 1280
rect 364198 800 364310 1280
rect 365380 0 365492 1280
rect 366562 800 366674 1280
rect 367744 800 367856 1280
rect 368926 0 369038 1280
rect 370108 800 370220 1280
rect 371290 800 371402 1280
rect 372472 0 372584 1280
rect 373654 800 373766 1280
rect 374836 800 374948 1280
rect 376018 0 376130 1280
rect 377200 800 377312 1280
rect 378382 800 378494 1280
rect 379564 0 379676 1280
rect 380746 800 380858 1280
rect 381928 800 382040 1280
rect 383110 0 383222 1280
rect 384292 800 384404 1280
rect 385474 800 385586 1280
rect 386656 0 386768 1280
rect 387838 800 387950 1280
rect 389020 800 389132 1280
rect 390202 0 390314 1280
rect 391384 800 391496 1280
rect 392566 800 392678 1280
rect 393748 0 393860 1280
rect 394930 800 395042 1280
rect 396112 800 396224 1280
rect 397294 0 397406 1280
rect 398476 800 398588 1280
rect 399658 800 399770 1280
rect 400840 0 400952 1280
rect 402022 800 402134 1280
rect 403204 800 403316 1280
rect 404386 0 404498 1280
rect 405568 800 405680 1280
rect 406750 800 406862 1280
rect 407932 0 408044 1280
rect 409114 800 409226 1280
rect 410296 800 410408 1280
rect 411478 0 411590 1280
rect 412660 800 412772 1280
rect 413842 800 413954 1280
rect 415024 0 415136 1280
rect 416206 800 416318 1280
rect 417388 800 417500 1280
rect 418570 0 418682 1280
rect 419752 800 419864 1280
rect 420934 800 421046 1280
rect 422116 0 422228 1280
rect 423298 800 423410 1280
rect 424480 800 424592 1280
rect 425662 0 425774 1280
rect 426844 800 426956 1280
rect 428026 800 428138 1280
rect 429205 1176 429325 2128
rect 432738 1280 432858 2128
rect 436289 1280 436406 2128
rect 439839 1280 439956 2128
rect 429208 0 429320 1176
rect 430390 800 430502 1280
rect 431572 800 431684 1280
rect 432738 1111 432866 1280
rect 432754 0 432866 1111
rect 433936 800 434048 1280
rect 435118 800 435230 1280
rect 436289 1014 436412 1280
rect 436300 0 436412 1014
rect 437482 800 437594 1280
rect 438664 800 438776 1280
rect 439839 981 439958 1280
rect 439846 0 439958 981
rect 441028 800 441140 1280
rect 442210 800 442322 1280
rect 443388 1014 443505 2128
rect 443392 0 443504 1014
rect 444574 800 444686 1280
rect 445756 800 445868 1280
rect 446938 1063 447055 2128
rect 448122 1280 448239 14561
rect 518034 14652 518114 605335
rect 560291 603833 560669 609925
rect 561257 609913 561263 610291
rect 561641 609913 561647 610291
rect 560282 603455 560291 603833
rect 560669 603455 560678 603833
rect 561263 602873 561641 609913
rect 561263 602486 561641 602495
rect 540027 598379 540281 598388
rect 540027 598116 540281 598125
rect 540098 524770 540218 598116
rect 563365 585567 563451 585576
rect 532586 522794 532670 522800
rect 450515 14496 450585 14500
rect 450488 14491 450605 14496
rect 450488 14421 450515 14491
rect 450585 14421 450605 14491
rect 450488 1280 450605 14421
rect 451699 14334 451769 14340
rect 451670 14331 451791 14334
rect 451670 14261 451699 14331
rect 451769 14261 451791 14331
rect 451670 1938 451791 14261
rect 518034 14240 518114 14572
rect 518194 522710 532586 522794
rect 518194 14488 518274 522710
rect 532586 522704 532670 522710
rect 532510 520290 532594 520296
rect 518194 14240 518274 14408
rect 518354 520206 532510 520290
rect 518354 14336 518434 520206
rect 532510 520200 532594 520206
rect 540184 512606 540304 513758
rect 540077 512597 540331 512606
rect 540077 512334 540331 512343
rect 530205 501603 530211 501689
rect 530297 501603 533953 501689
rect 534039 501603 534048 501689
rect 563365 501684 563451 585481
rect 571878 584670 571948 585410
rect 563365 501608 563370 501684
rect 563446 501608 563451 501684
rect 563365 501603 563451 501608
rect 565274 584590 571948 584670
rect 563370 501599 563446 501603
rect 530697 501247 530783 501253
rect 530783 501161 533965 501247
rect 534051 501161 534060 501247
rect 530697 501155 530783 501161
rect 541397 488631 542206 488831
rect 542406 488631 542415 488831
rect 544533 488260 544619 488266
rect 544619 488174 550031 488260
rect 550117 488174 550126 488260
rect 544533 488168 544619 488174
rect 542134 481594 542186 481600
rect 542134 481536 542186 481542
rect 541946 480616 541952 480668
rect 542004 480616 542010 480668
rect 541960 479524 541996 480616
rect 523634 479488 541996 479524
rect 523474 388631 523554 388634
rect 520412 388626 523554 388631
rect 520408 388500 520417 388626
rect 520543 388500 523554 388626
rect 520412 388495 523554 388500
rect 520134 387923 523334 387928
rect 520130 387797 520139 387923
rect 520265 387797 523334 387923
rect 520134 387792 523334 387797
rect 519109 386264 519235 386268
rect 523094 386264 523174 386268
rect 519104 386259 523174 386264
rect 519104 386133 519109 386259
rect 519235 386133 523174 386259
rect 519104 386128 523174 386133
rect 519109 386124 519235 386128
rect 520091 385247 520217 385251
rect 522934 385247 523014 385252
rect 520086 385242 523014 385247
rect 520086 385116 520091 385242
rect 520217 385116 523014 385242
rect 520086 385111 523014 385116
rect 520091 385107 520217 385111
rect 520796 383269 520860 383273
rect 522774 383269 522854 383270
rect 520791 383264 522854 383269
rect 520791 383200 520796 383264
rect 520860 383200 522854 383264
rect 520791 383195 522854 383200
rect 520796 383191 520860 383195
rect 521200 380963 521256 380970
rect 522554 380963 522634 380964
rect 521198 380961 522634 380963
rect 521198 380905 521200 380961
rect 521256 380905 522634 380961
rect 521198 380903 522634 380905
rect 521200 380896 521256 380903
rect 519146 378844 519202 378851
rect 522394 378844 522474 378848
rect 519144 378842 522474 378844
rect 519144 378786 519146 378842
rect 519202 378786 522474 378842
rect 519144 378784 522474 378786
rect 519146 378777 519202 378784
rect 519085 378591 522314 378596
rect 519081 378507 519090 378591
rect 519174 378507 522314 378591
rect 519085 378502 522314 378507
rect 519150 378368 519234 378372
rect 522074 378368 522154 378370
rect 519145 378363 522154 378368
rect 519145 378279 519150 378363
rect 519234 378279 522154 378363
rect 519145 378274 522154 378279
rect 519150 378270 519234 378274
rect 519290 378086 519374 378090
rect 519285 378081 521934 378086
rect 519285 377997 519290 378081
rect 519374 377997 521934 378081
rect 519285 377992 521934 377997
rect 519290 377988 519374 377992
rect 521694 375546 521774 375548
rect 518978 375466 518984 375546
rect 519064 375466 521774 375546
rect 521534 372934 521614 372936
rect 520740 372854 520746 372934
rect 520826 372854 521614 372934
rect 521374 367944 521454 367946
rect 520834 367864 520840 367944
rect 520920 367864 521454 367944
rect 521154 349350 521234 349384
rect 520994 349040 521074 349068
rect 520834 348700 520914 348730
rect 520674 348348 520754 348380
rect 520454 348062 520534 348128
rect 520294 347814 520374 347878
rect 520134 347548 520214 347600
rect 519974 347284 520054 347338
rect 519754 313970 519834 314022
rect 519594 313516 519674 313568
rect 519434 313164 519514 313198
rect 519274 312776 519354 312872
rect 519054 312230 519134 312308
rect 518894 311660 518974 311746
rect 518734 311230 518814 311342
rect 518354 14240 518434 14256
rect 518574 310692 518654 310820
rect 454049 14191 454139 14200
rect 451672 1280 451789 1938
rect 454049 1280 454139 14101
rect 518574 14174 518654 310612
rect 455233 14025 455323 14034
rect 455233 1280 455323 13935
rect 457581 13857 457671 13866
rect 457581 1280 457671 13767
rect 458765 13699 458855 13708
rect 458765 1280 458855 13609
rect 518574 13570 518654 14094
rect 518734 14022 518814 311150
rect 518734 13570 518814 13942
rect 518894 13858 518974 311580
rect 518894 13570 518974 13778
rect 519054 13696 519134 312150
rect 519054 13570 519134 13616
rect 461132 13539 461222 13548
rect 461132 1280 461222 13449
rect 519274 13528 519354 312696
rect 462316 13381 462406 13390
rect 462316 1280 462406 13291
rect 464676 13226 464760 13235
rect 464676 1280 464760 13142
rect 465851 12976 465860 13060
rect 465944 12976 465953 13060
rect 465860 1280 465944 12976
rect 519274 12922 519354 13448
rect 519434 13374 519514 313084
rect 519434 12922 519514 13294
rect 519594 13216 519674 313436
rect 519594 12922 519674 13136
rect 519754 13056 519834 313890
rect 519754 12922 519834 12976
rect 468227 12894 468311 12903
rect 468227 1280 468311 12810
rect 519974 12898 520054 347204
rect 469411 12738 469495 12747
rect 469411 1280 469495 12654
rect 471768 12574 471852 12583
rect 471768 1280 471852 12490
rect 472952 12414 473036 12423
rect 472952 1280 473036 12330
rect 519974 12274 520054 12818
rect 520134 12738 520214 347468
rect 520134 12274 520214 12658
rect 520294 12578 520374 347734
rect 520294 12274 520374 12498
rect 520454 12418 520534 347982
rect 520454 12274 520534 12338
rect 475319 12264 475403 12273
rect 475319 1280 475403 12180
rect 520674 12256 520754 348268
rect 476503 12100 476587 12109
rect 476503 1280 476587 12016
rect 478869 11940 478953 11949
rect 478869 1280 478953 11856
rect 480053 11782 480137 11791
rect 480053 1280 480137 11698
rect 520674 11664 520754 12176
rect 520834 12098 520914 348620
rect 520834 11664 520914 12018
rect 520994 11936 521074 348960
rect 520994 11664 521074 11856
rect 521154 11776 521234 349270
rect 521154 11664 521234 11696
rect 482415 11621 482490 11630
rect 482415 1280 482490 11546
rect 521374 11614 521454 367864
rect 483599 11455 483674 11464
rect 483599 1280 483674 11380
rect 485956 11299 486031 11308
rect 485956 1280 486031 11224
rect 487140 11139 487215 11148
rect 487140 1280 487215 11064
rect 521374 10992 521454 11534
rect 521534 11458 521614 372854
rect 521534 10992 521614 11378
rect 521694 11288 521774 375466
rect 521694 10992 521774 11208
rect 521854 11136 521934 377992
rect 521854 10992 521934 11056
rect 489478 10973 489553 10982
rect 489478 1280 489553 10898
rect 522074 10974 522154 378274
rect 490662 10817 490737 10826
rect 490662 1280 490737 10742
rect 493048 10655 493123 10664
rect 493048 1280 493123 10580
rect 494232 10499 494307 10508
rect 494232 1280 494307 10424
rect 522074 10370 522154 10894
rect 522234 10810 522314 378502
rect 522234 10370 522314 10730
rect 522394 10652 522474 378784
rect 522394 10370 522474 10572
rect 522554 10494 522634 380903
rect 522554 10370 522634 10414
rect 496589 10327 496664 10336
rect 496589 1280 496664 10252
rect 522774 10332 522854 383195
rect 497773 10171 497848 10180
rect 497773 1280 497848 10096
rect 500140 10015 500215 10024
rect 500140 1280 500215 9940
rect 501324 9851 501399 9860
rect 501324 1280 501399 9776
rect 522774 9710 522854 10252
rect 522934 10178 523014 385111
rect 522934 9710 523014 10098
rect 523094 10026 523174 386128
rect 523094 9710 523174 9946
rect 523254 9852 523334 387792
rect 523254 9710 523334 9772
rect 503689 9684 503749 9693
rect 503689 9615 503749 9624
rect 523474 9690 523554 388495
rect 503690 1280 503748 9615
rect 504873 9524 504933 9533
rect 504873 9455 504933 9464
rect 504874 1280 504932 9455
rect 507249 9368 507309 9377
rect 507249 9299 507309 9308
rect 507250 1280 507308 9299
rect 508433 9216 508493 9225
rect 508433 9147 508493 9156
rect 508434 1280 508492 9147
rect 523474 9074 523554 9610
rect 523634 9538 523714 479488
rect 542142 479406 542178 481536
rect 523634 9074 523714 9458
rect 523794 479370 542178 479406
rect 523794 9370 523874 479370
rect 553602 376077 556571 376083
rect 549547 373108 549556 376077
rect 552525 373108 553602 376077
rect 553602 373102 556571 373108
rect 563162 260786 563802 260862
rect 563878 260786 563887 260862
rect 524985 256303 524994 256611
rect 525302 256303 527559 256611
rect 563238 256438 563738 256514
rect 563814 256438 563823 256514
rect 563596 255774 564753 256071
rect 562858 255696 564753 255774
rect 562858 255399 563971 255696
rect 563228 254912 563752 254988
rect 563828 254912 563837 254988
rect 524547 253131 524556 253331
rect 524756 253131 527556 253331
rect 524670 252435 524679 252974
rect 525218 252435 527890 252974
rect 564378 244544 564753 255696
rect 562630 244169 562639 244544
rect 563014 244169 564753 244544
rect 552198 170461 552369 170467
rect 552369 170290 558218 170461
rect 558389 170290 558398 170461
rect 552198 170284 552369 170290
rect 523794 9074 523874 9290
rect 523954 152725 535546 152728
rect 523954 152667 535443 152725
rect 535501 152667 535546 152725
rect 523954 152648 535546 152667
rect 523954 9216 524034 152648
rect 523954 9074 524034 9136
rect 524174 152493 537146 152508
rect 524174 152435 537071 152493
rect 537129 152435 537146 152493
rect 524174 152428 537146 152435
rect 510800 9046 510860 9055
rect 510800 8977 510860 8986
rect 524174 9054 524254 152428
rect 510801 1280 510859 8977
rect 511984 8886 512044 8895
rect 511984 8817 512044 8826
rect 511985 1280 512043 8817
rect 514324 8730 514400 8739
rect 514324 1280 514400 8654
rect 515508 8570 515584 8579
rect 515508 1280 515584 8494
rect 524174 8440 524254 8974
rect 524334 152343 538794 152348
rect 524334 152285 538699 152343
rect 538757 152285 538794 152343
rect 524334 152268 538794 152285
rect 524334 8896 524414 152268
rect 524334 8440 524414 8816
rect 524494 152179 540428 152188
rect 524494 152121 540327 152179
rect 540385 152121 540428 152179
rect 524494 152108 540428 152121
rect 524494 8738 524574 152108
rect 524494 8440 524574 8658
rect 524654 152025 542068 152028
rect 524654 151967 541955 152025
rect 542013 151967 542068 152025
rect 524654 151948 542068 151967
rect 524654 8570 524734 151948
rect 524654 8440 524734 8490
rect 524874 151787 543696 151808
rect 524874 151729 543583 151787
rect 543641 151729 543696 151787
rect 524874 151728 543696 151729
rect 517874 8414 517950 8423
rect 517874 1280 517950 8338
rect 524874 8414 524954 151728
rect 519058 8254 519134 8263
rect 519058 1280 519134 8178
rect 521425 8090 521501 8099
rect 521425 1280 521501 8014
rect 522609 7930 522685 7939
rect 522609 1280 522685 7854
rect 524874 7832 524954 8334
rect 525034 151633 545330 151648
rect 525034 151575 545211 151633
rect 545269 151575 545330 151633
rect 525034 151568 545330 151575
rect 525034 8260 525114 151568
rect 525034 7832 525114 8180
rect 525194 151475 546928 151488
rect 525194 151417 546839 151475
rect 546897 151417 546928 151475
rect 525194 151408 546928 151417
rect 548994 151435 549287 155046
rect 525194 8096 525274 151408
rect 548994 151133 549287 151142
rect 549439 150748 549818 154995
rect 549439 150360 549818 150369
rect 557518 73522 558751 73648
rect 558877 73522 558886 73648
rect 536989 56451 536995 56509
rect 537053 56451 537059 56509
rect 536995 53783 537053 56451
rect 538617 56327 538623 56385
rect 538681 56327 538687 56385
rect 540245 56349 540251 56407
rect 540309 56349 540315 56407
rect 538623 53973 538681 56327
rect 540251 55739 540309 56349
rect 541873 56331 541879 56389
rect 541937 56331 541943 56389
rect 540010 55738 540309 55739
rect 539734 55681 540309 55738
rect 539574 53973 539654 53974
rect 538623 53915 539654 53973
rect 536995 53725 539435 53783
rect 525194 7832 525274 8016
rect 539354 7940 539434 53725
rect 539354 7804 539434 7860
rect 524976 7772 525052 7781
rect 524976 1280 525052 7696
rect 539574 7778 539654 53915
rect 526160 7616 526236 7625
rect 526160 1280 526236 7540
rect 528508 7458 528584 7467
rect 528508 1280 528584 7382
rect 529692 7302 529768 7311
rect 529692 1280 529768 7226
rect 539574 7170 539654 7698
rect 539734 7624 539814 55681
rect 541879 55534 541937 56331
rect 543501 56267 543507 56325
rect 543565 56267 543571 56325
rect 539734 7170 539814 7544
rect 539894 55477 541937 55534
rect 539894 55454 541936 55477
rect 539894 7466 539974 55454
rect 543507 55336 543565 56267
rect 546757 56239 546763 56297
rect 546821 56239 546827 56297
rect 545135 56197 545193 56203
rect 539894 7170 539974 7386
rect 540054 55256 543566 55336
rect 540054 7294 540134 55256
rect 545135 55108 545193 56139
rect 540054 7170 540134 7214
rect 540274 55028 545194 55108
rect 532049 7142 532125 7151
rect 532049 1280 532125 7066
rect 540274 7142 540354 55028
rect 546763 54904 546821 56239
rect 548385 56195 548391 56253
rect 548449 56195 548455 56253
rect 549825 56202 549831 56254
rect 549883 56202 549889 56254
rect 533233 6972 533309 6981
rect 533233 1280 533309 6896
rect 535609 6824 535685 6833
rect 535609 1280 535685 6748
rect 536793 6648 536869 6657
rect 536793 1280 536869 6572
rect 540274 6546 540354 7062
rect 540434 54824 546822 54904
rect 540434 6976 540514 54824
rect 548391 54682 548449 56195
rect 540434 6546 540514 6896
rect 540594 54603 548449 54682
rect 549839 54644 549875 56202
rect 550546 55249 550839 56731
rect 550546 54947 550839 54956
rect 550991 54732 551370 56817
rect 540594 54602 548446 54603
rect 540594 6816 540674 54602
rect 549798 54456 549878 54644
rect 540594 6546 540674 6736
rect 540754 54376 549878 54456
rect 540754 6662 540834 54376
rect 550991 54344 551370 54353
rect 540754 6546 540834 6582
rect 539150 6496 539226 6526
rect 550274 6512 550354 6546
rect 550434 6512 550514 6546
rect 550594 6512 550674 6546
rect 550754 6512 550834 6546
rect 539150 1280 539226 6420
rect 565274 6498 565354 584590
rect 572018 584510 572088 585410
rect 540334 6324 540410 6370
rect 540334 1280 540410 6248
rect 542706 6172 542783 6194
rect 541522 1280 541599 1340
rect 542706 1280 542783 6095
rect 543890 6012 543967 6040
rect 543890 1280 543967 5935
rect 565274 5886 565354 6418
rect 565434 584430 572088 584510
rect 565434 6344 565514 584430
rect 572158 584350 572228 585410
rect 565434 5886 565514 6264
rect 565594 584270 572228 584350
rect 565594 6180 565674 584270
rect 572298 584190 572368 585410
rect 565594 5886 565674 6100
rect 565754 584110 572368 584190
rect 565754 6014 565834 584110
rect 571878 503870 571948 504610
rect 565754 5886 565834 5934
rect 566274 503790 571948 503870
rect 546251 5860 546328 5880
rect 545067 1280 545144 1314
rect 546251 1280 546328 5783
rect 566274 5854 566354 503790
rect 572018 503710 572088 504610
rect 547435 5700 547512 5718
rect 547435 1280 547512 5623
rect 549788 5528 549865 5558
rect 548604 1280 548681 1332
rect 549788 1280 549865 5451
rect 550972 5372 551049 5386
rect 550972 1280 551049 5295
rect 566274 5264 566354 5774
rect 566434 503630 572088 503710
rect 566434 5700 566514 503630
rect 572158 503550 572228 504610
rect 566434 5264 566514 5620
rect 566594 503470 572228 503550
rect 566594 5542 566674 503470
rect 572298 503390 572368 504610
rect 566594 5264 566674 5462
rect 566754 503310 572368 503390
rect 566754 5380 566834 503310
rect 571878 487470 571948 488210
rect 566754 5264 566834 5300
rect 567274 487390 571948 487470
rect 553346 5218 553423 5236
rect 552162 1280 552239 1302
rect 553346 1280 553423 5141
rect 567274 5216 567354 487390
rect 572018 487310 572088 488210
rect 554530 5046 554607 5072
rect 554530 1280 554607 4969
rect 556886 4894 556970 4926
rect 556886 1280 556970 4810
rect 558070 4734 558154 4754
rect 558070 1280 558154 4650
rect 560405 4571 560525 4612
rect 567274 4604 567354 5136
rect 567434 487230 572088 487310
rect 567434 5060 567514 487230
rect 572158 487150 572228 488210
rect 567434 4604 567514 4980
rect 567594 487070 572228 487150
rect 567594 4902 567674 487070
rect 572298 486990 572368 488210
rect 567594 4604 567674 4822
rect 567754 486910 572368 486990
rect 567754 4732 567834 486910
rect 571878 471070 571948 471810
rect 567754 4604 567834 4652
rect 568274 470990 571948 471070
rect 560405 4501 560425 4571
rect 560495 4501 560525 4571
rect 560405 1445 560525 4501
rect 568274 4574 568354 470990
rect 572018 470910 572088 471810
rect 561589 4411 561709 4450
rect 561589 4341 561625 4411
rect 561695 4341 561709 4411
rect 448120 1063 448239 1280
rect 446938 0 447050 1063
rect 448120 800 448232 1063
rect 449302 800 449414 1280
rect 450484 1096 450605 1280
rect 451666 1096 451789 1280
rect 450484 0 450596 1096
rect 451666 800 451778 1096
rect 452848 800 452960 1280
rect 454019 1122 454142 1280
rect 454030 0 454142 1122
rect 455212 800 455324 1280
rect 456394 800 456506 1280
rect 457576 1190 457696 1280
rect 455233 0 455323 800
rect 457576 0 457688 1190
rect 458758 800 458870 1280
rect 459940 800 460052 1280
rect 461112 1086 461234 1280
rect 458765 0 458855 800
rect 461122 0 461234 1086
rect 462304 800 462416 1280
rect 463486 800 463598 1280
rect 464668 1094 464787 1280
rect 462316 0 462406 800
rect 464668 0 464780 1094
rect 465850 800 465962 1280
rect 467032 800 467144 1280
rect 468212 1163 468329 1280
rect 465860 0 465944 800
rect 468214 0 468326 1163
rect 469396 800 469508 1280
rect 470578 800 470690 1280
rect 471754 1147 471872 1280
rect 469411 0 469495 800
rect 471760 0 471872 1147
rect 472942 800 473054 1280
rect 474124 800 474236 1280
rect 475296 1117 475418 1280
rect 472952 0 473036 800
rect 475306 0 475418 1117
rect 476488 800 476600 1280
rect 477670 800 477782 1280
rect 476503 0 476587 800
rect 478852 0 478964 1280
rect 480034 800 480146 1280
rect 481216 800 481328 1280
rect 480053 0 480137 800
rect 482398 0 482510 1280
rect 483580 800 483692 1280
rect 484762 800 484874 1280
rect 483599 0 483674 800
rect 485944 0 486056 1280
rect 487126 800 487238 1280
rect 488308 800 488420 1280
rect 489478 1124 489602 1280
rect 490662 1124 490784 1280
rect 487140 0 487215 800
rect 489490 0 489602 1124
rect 490672 800 490784 1124
rect 491854 800 491966 1280
rect 493036 0 493148 1280
rect 494218 800 494330 1280
rect 495400 800 495512 1280
rect 494232 0 494307 800
rect 496582 0 496694 1280
rect 497764 800 497876 1280
rect 498946 800 499058 1280
rect 497773 0 497848 800
rect 500128 0 500240 1280
rect 501310 800 501422 1280
rect 502492 800 502604 1280
rect 501324 0 501399 800
rect 503674 0 503786 1280
rect 504856 800 504968 1280
rect 506038 800 506150 1280
rect 504874 0 504932 800
rect 507220 0 507332 1280
rect 508402 800 508514 1280
rect 509584 800 509696 1280
rect 508434 0 508492 800
rect 510766 0 510878 1280
rect 511948 800 512060 1280
rect 513130 800 513242 1280
rect 511985 0 512043 800
rect 514312 0 514424 1280
rect 515494 800 515606 1280
rect 516676 800 516788 1280
rect 515508 0 515584 800
rect 517858 0 517970 1280
rect 519040 800 519152 1280
rect 520222 800 520334 1280
rect 519058 0 519134 800
rect 521404 0 521516 1280
rect 522586 800 522698 1280
rect 523768 800 523880 1280
rect 522609 0 522685 800
rect 524950 0 525062 1280
rect 526132 800 526244 1280
rect 527314 800 527426 1280
rect 526160 0 526236 800
rect 528496 0 528608 1280
rect 529678 800 529790 1280
rect 530860 800 530972 1280
rect 529692 0 529768 800
rect 532042 0 532154 1280
rect 533224 800 533336 1280
rect 534406 800 534518 1280
rect 533233 0 533309 800
rect 535588 0 535700 1280
rect 536770 800 536882 1280
rect 537952 800 538064 1280
rect 536793 0 536869 800
rect 539134 0 539246 1280
rect 540316 800 540428 1280
rect 540334 0 540410 800
rect 541498 0 541610 1280
rect 542680 800 542792 1280
rect 543862 800 543974 1280
rect 542706 0 542783 800
rect 543890 0 543967 800
rect 545044 0 545156 1280
rect 546226 800 546338 1280
rect 547408 800 547520 1280
rect 546251 0 546328 800
rect 547435 0 547512 800
rect 548590 0 548702 1280
rect 549772 800 549884 1280
rect 550954 800 551066 1280
rect 549788 0 549865 800
rect 550972 0 551049 800
rect 552136 0 552248 1280
rect 553318 800 553430 1280
rect 554500 800 554612 1280
rect 555682 800 555794 1280
rect 553346 0 553423 800
rect 554530 0 554607 800
rect 556864 0 556976 1280
rect 558046 800 558158 1280
rect 559228 800 559340 1280
rect 558070 0 558154 800
rect 560410 0 560522 1445
rect 561589 1174 561709 4341
rect 563980 4262 564056 4284
rect 563980 1280 564056 4186
rect 565164 4102 565240 4142
rect 565164 1280 565240 4026
rect 567527 3941 567605 3951
rect 568274 3946 568354 4494
rect 568434 470830 572088 470910
rect 568434 4408 568514 470830
rect 572158 470750 572228 471810
rect 568434 3946 568514 4328
rect 568594 470670 572228 470750
rect 568594 4250 568674 470670
rect 572298 470590 572368 471810
rect 568594 3946 568674 4170
rect 568754 470510 572368 470590
rect 568754 4092 568834 470510
rect 577992 360764 577998 363733
rect 580967 360764 580973 363733
rect 577998 356751 580967 360764
rect 577998 353773 580967 353782
rect 571878 309670 571948 310410
rect 568754 3946 568834 4012
rect 569274 309590 571948 309670
rect 567527 1280 567605 3863
rect 569274 3924 569354 309590
rect 572018 309510 572088 310410
rect 568711 3773 568789 3782
rect 568711 1280 568789 3695
rect 569274 3334 569354 3844
rect 569434 309430 572088 309510
rect 569434 3772 569514 309430
rect 572158 309350 572228 310410
rect 569434 3334 569514 3692
rect 569594 309270 572228 309350
rect 569594 3612 569674 309270
rect 572298 309190 572368 310410
rect 569594 3334 569674 3532
rect 569754 309110 572368 309190
rect 569754 3454 569834 309110
rect 571878 270070 571948 270722
rect 569754 3334 569834 3374
rect 570274 269990 571948 270070
rect 570274 3298 570354 269990
rect 572018 269910 572088 270722
rect 570274 2620 570354 3218
rect 570434 269830 572088 269910
rect 570434 3136 570514 269830
rect 572158 269750 572228 270722
rect 570434 2620 570514 3056
rect 570594 269670 572228 269750
rect 570594 2976 570674 269670
rect 572298 269590 572368 270722
rect 570594 2620 570674 2896
rect 570754 269510 572368 269590
rect 570754 2808 570834 269510
rect 570754 2620 570834 2728
rect 571050 3615 571128 3657
rect 571050 1280 571128 3537
rect 572234 3461 572312 3491
rect 572234 1280 572312 3383
rect 574610 3295 574688 3349
rect 574610 1280 574688 3217
rect 575794 3139 575872 3181
rect 575794 1280 575872 3061
rect 578154 2977 578232 2997
rect 578154 1280 578232 2899
rect 579338 2815 579416 2855
rect 579338 1280 579416 2737
rect 561592 800 561704 1174
rect 562774 800 562886 1280
rect 563956 0 564068 1280
rect 565138 800 565250 1280
rect 566320 800 566432 1280
rect 565164 0 565240 800
rect 567502 0 567614 1280
rect 568684 800 568796 1280
rect 569866 800 569978 1280
rect 568711 0 568789 800
rect 571048 0 571160 1280
rect 572230 800 572342 1280
rect 573412 800 573524 1280
rect 574594 800 574706 1280
rect 575776 800 575888 1280
rect 576958 800 577070 1280
rect 578140 800 578252 1280
rect 579322 800 579434 1280
rect 580504 800 580616 1280
rect 581686 800 581798 1280
rect 582868 800 582980 1280
rect 584050 800 584162 1280
rect 572234 0 572312 800
rect 575794 0 575872 800
rect 579338 0 579416 800
<< via2 >>
rect 138173 656216 139419 657462
rect 445405 656216 446651 657462
rect 130007 653816 131253 655062
rect 453593 653816 454839 655062
rect 12714 2009 12784 2079
rect 12854 2177 12924 2247
rect 12994 2337 13064 2407
rect 13734 2653 13804 2723
rect 13894 2813 13964 2883
rect 14054 2973 14124 3043
rect 14734 3293 14804 3363
rect 14894 3449 14964 3519
rect 15054 3615 15124 3685
rect 15734 3929 15804 3999
rect 15894 4097 15964 4167
rect 16054 4257 16124 4327
rect 16734 4567 16804 4637
rect 16894 4729 16964 4799
rect 17054 4893 17124 4963
rect 17734 5211 17804 5281
rect 17894 5373 17964 5443
rect 18054 5537 18124 5607
rect 18734 5849 18804 5919
rect 18894 6013 18964 6083
rect 19054 6177 19124 6247
rect 19734 6493 19804 6563
rect 19894 6655 19964 6725
rect 20054 6815 20124 6885
rect 20734 7133 20804 7203
rect 20894 7291 20964 7361
rect 21054 7451 21124 7521
rect 21734 7775 21804 7845
rect 21894 7935 21964 8005
rect 22054 8097 22124 8167
rect 32420 496192 32488 496260
rect 70696 496202 70780 496286
rect 30866 494838 31406 495378
rect 32714 494100 32774 494160
rect 31040 492746 31580 493286
rect 32716 491588 32772 491644
rect 32425 491437 32483 491495
rect 34415 468421 34669 468675
rect 28647 437183 28901 437437
rect 33711 467715 33965 467969
rect 32303 424515 32557 424769
rect 55450 426023 55650 426223
rect 55426 424701 55626 424901
rect 55428 424396 55628 424596
rect 37908 412714 38108 412914
rect 32967 381315 33221 381569
rect 23112 350708 23212 350808
rect 40087 334472 40593 334978
rect 40079 333578 40561 334060
rect 38766 331899 38866 331999
rect 24332 331339 24432 331439
rect 23124 307420 23224 307520
rect 40653 283675 42243 285265
rect 45657 276361 47247 277951
rect 39312 222735 39964 223387
rect 61931 223542 62593 224204
rect 45947 222730 46609 223392
rect 61877 222730 62539 223392
rect 44023 132506 45134 133617
rect 50123 131168 50501 131546
rect 42543 130699 42645 130801
rect 50097 128787 50475 129165
rect 44572 126745 45683 127856
rect 41188 58143 42568 59523
rect 42439 57188 42509 57258
rect 42429 9441 42531 9543
rect 42745 57008 42815 57078
rect 42743 9045 42845 9147
rect 70734 8413 70804 8483
rect 70894 8573 70964 8643
rect 71054 8733 71124 8803
rect 71434 9051 71504 9121
rect 71594 9215 71664 9285
rect 71754 9375 71824 9445
rect 72134 9695 72204 9765
rect 72294 9855 72364 9925
rect 72454 10015 72524 10085
rect 72834 10335 72904 10405
rect 72994 10495 73064 10565
rect 73154 10653 73224 10723
rect 73534 10977 73604 11047
rect 73694 11131 73764 11201
rect 73854 11293 73924 11363
rect 74234 11611 74304 11681
rect 74394 11775 74464 11845
rect 74554 11933 74624 12003
rect 74934 12255 75004 12325
rect 75094 12411 75164 12481
rect 75254 12573 75324 12643
rect 75634 12893 75704 12963
rect 75794 13051 75864 13121
rect 75954 13213 76024 13283
rect 126893 591344 127014 591465
rect 138287 566216 139533 567462
rect 130007 563816 131253 565062
rect 130498 520258 130794 520554
rect 138463 519191 138773 519501
rect 138401 476216 139647 477462
rect 130159 473816 131405 475062
rect 138267 386216 139513 387462
rect 130159 383816 131405 385062
rect 138115 296216 139361 297462
rect 129929 293816 131175 295062
rect 138191 206216 139437 207462
rect 130159 203816 131405 205062
rect 138173 116216 139419 117462
rect 130007 113816 131253 115062
rect 76114 13377 76184 13447
rect 253096 13374 253167 13445
rect 251904 13214 251975 13285
rect 249554 13054 249625 13125
rect 248370 12894 248441 12965
rect 75414 12733 75484 12803
rect 246011 12721 246101 12811
rect 244827 12561 244917 12651
rect 242475 12407 242565 12497
rect 241291 12245 241381 12335
rect 74714 12091 74784 12161
rect 238927 12083 239017 12173
rect 237743 11921 237833 12011
rect 235362 11754 235462 11854
rect 234178 11596 234278 11696
rect 74014 11453 74084 11523
rect 231814 11442 231914 11542
rect 230630 11284 230730 11384
rect 228288 11124 228388 11224
rect 227104 10960 227204 11060
rect 73314 10813 73384 10883
rect 224740 10800 224840 10900
rect 223556 10642 223656 10742
rect 221202 10484 221302 10584
rect 220018 10322 220118 10422
rect 72614 10173 72684 10243
rect 217658 10174 217729 10245
rect 216476 10014 216547 10085
rect 214129 9851 214198 9920
rect 212945 9689 213014 9758
rect 71914 9537 71984 9607
rect 210577 9527 210646 9596
rect 209393 9369 209462 9438
rect 207019 9223 207088 9292
rect 205835 9065 205904 9134
rect 71214 8893 71284 8963
rect 203478 8900 203538 8960
rect 202294 8742 202354 8802
rect 199920 8571 200010 8661
rect 198736 8401 198826 8491
rect 22214 8253 22284 8323
rect 196359 8249 196449 8339
rect 195175 8083 195265 8173
rect 192827 7921 192897 7991
rect 191643 7779 191713 7849
rect 21214 7613 21284 7683
rect 189287 7613 189368 7694
rect 188103 7439 188184 7520
rect 185747 7291 185828 7372
rect 184563 7137 184644 7218
rect 20214 6975 20284 7045
rect 182183 6969 182264 7050
rect 180999 6815 181080 6896
rect 178632 6651 178713 6732
rect 177448 6493 177529 6574
rect 19214 6333 19284 6403
rect 175093 6327 175174 6408
rect 173909 6167 173990 6248
rect 171566 6013 171647 6094
rect 170382 5849 170463 5930
rect 18214 5693 18284 5763
rect 168002 5687 168083 5768
rect 166818 5527 166899 5608
rect 164457 5365 164538 5446
rect 163273 5221 163354 5302
rect 17214 5053 17284 5123
rect 160918 5043 160999 5124
rect 159734 4875 159815 4956
rect 157360 4725 157441 4806
rect 156176 4571 156257 4652
rect 16214 4419 16284 4489
rect 153808 4407 153889 4488
rect 152624 4253 152705 4334
rect 150282 4089 150363 4170
rect 149098 3927 149179 4008
rect 15214 3771 15284 3841
rect 146724 3771 146805 3852
rect 145540 3613 145621 3694
rect 143191 3453 143272 3534
rect 142007 3287 142088 3368
rect 14214 3129 14284 3199
rect 139633 3135 139714 3216
rect 138449 2969 138530 3050
rect 136088 2819 136169 2900
rect 134904 2647 134985 2728
rect 13134 2493 13204 2563
rect 132555 2481 132636 2562
rect 131371 2325 131452 2406
rect 129002 2179 129083 2260
rect 127818 2007 127899 2088
rect 280296 9876 280356 9936
rect 276749 9700 276809 9760
rect 273201 9550 273261 9610
rect 282707 10484 282767 10544
rect 294486 10508 294546 10568
rect 282427 10346 282487 10406
rect 290938 10350 290998 10410
rect 282147 10168 282207 10228
rect 287391 10192 287451 10252
rect 281867 10006 281927 10066
rect 283843 10042 283903 10102
rect 281587 9852 281647 9912
rect 281307 9690 281367 9750
rect 281027 9528 281087 9588
rect 298033 9380 298093 9440
rect 538251 613613 540245 615607
rect 583269 611592 583343 611666
rect 541059 606980 543053 608974
rect 454034 592807 454330 593103
rect 445481 566216 446727 567462
rect 453515 563816 454761 565062
rect 303962 9382 304022 9442
rect 301569 9222 301629 9282
rect 445841 494877 446151 495187
rect 454080 483040 454376 483336
rect 445367 476216 446613 477462
rect 453439 473816 454685 475062
rect 304242 9212 304302 9272
rect 517544 388495 517680 388631
rect 517556 387792 517692 387928
rect 445481 386216 446727 387462
rect 517688 386128 517824 386264
rect 517526 385111 517662 385247
rect 453515 383816 454761 385062
rect 516805 383195 516879 383269
rect 451716 382153 451776 382213
rect 438563 381198 438742 381377
rect 304522 9058 304582 9118
rect 439337 381257 439555 381475
rect 439833 381255 439963 381385
rect 441444 381051 442145 381752
rect 442634 381019 443287 381672
rect 451236 381134 451372 381270
rect 506922 380903 506982 380963
rect 516870 378784 516930 378844
rect 516821 378502 516915 378596
rect 516881 378274 516975 378368
rect 516953 377992 517047 378086
rect 461915 377649 462017 377751
rect 461195 377283 461297 377385
rect 505921 376821 506251 377151
rect 450424 376009 450836 376421
rect 449325 374677 449759 375111
rect 490958 349242 491094 349378
rect 490906 348922 491042 349058
rect 490890 348584 491026 348720
rect 490958 348230 491094 348366
rect 490822 347960 490958 348096
rect 490822 347706 490958 347842
rect 490890 347436 491026 347572
rect 490940 347166 491076 347302
rect 445367 296216 446613 297462
rect 453707 293816 454953 295062
rect 304802 8896 304862 8956
rect 445597 206216 446843 207462
rect 453325 203816 454571 205062
rect 305082 8718 305142 8778
rect 445481 116216 446727 117462
rect 453593 113816 454839 115062
rect 305362 8572 305422 8632
rect 448122 14561 448239 14678
rect 305642 8426 305702 8486
rect 306122 9068 306182 9128
rect 308682 8902 308742 8962
rect 312210 8750 312270 8810
rect 315770 8600 315830 8660
rect 319309 8424 319369 8484
rect 560291 603455 560669 603833
rect 561263 602495 561641 602873
rect 540027 598125 540281 598379
rect 563365 585481 563451 585567
rect 518034 14572 518114 14652
rect 450515 14421 450585 14491
rect 451699 14261 451769 14331
rect 518194 14408 518274 14488
rect 540077 512343 540331 512597
rect 533953 501603 534039 501689
rect 563370 501608 563446 501684
rect 533965 501161 534051 501247
rect 542206 488631 542406 488831
rect 550031 488174 550117 488260
rect 520417 388500 520543 388626
rect 520139 387797 520265 387923
rect 519109 386133 519235 386259
rect 520091 385116 520217 385242
rect 520796 383200 520860 383264
rect 521200 380905 521256 380961
rect 519146 378786 519202 378842
rect 519090 378507 519174 378591
rect 519150 378279 519234 378363
rect 519290 377997 519374 378081
rect 521154 349270 521234 349350
rect 520994 348960 521074 349040
rect 520834 348620 520914 348700
rect 520674 348268 520754 348348
rect 520454 347982 520534 348062
rect 520294 347734 520374 347814
rect 520134 347468 520214 347548
rect 519974 347204 520054 347284
rect 518354 14256 518434 14336
rect 454049 14101 454139 14191
rect 518574 14094 518654 14174
rect 455233 13935 455323 14025
rect 457581 13767 457671 13857
rect 458765 13609 458855 13699
rect 518734 13942 518814 14022
rect 518894 13778 518974 13858
rect 519054 13616 519134 13696
rect 461132 13449 461222 13539
rect 519274 13448 519354 13528
rect 462316 13291 462406 13381
rect 464676 13142 464760 13226
rect 465860 12976 465944 13060
rect 519434 13294 519514 13374
rect 519594 13136 519674 13216
rect 519754 12976 519834 13056
rect 468227 12810 468311 12894
rect 519974 12818 520054 12898
rect 469411 12654 469495 12738
rect 471768 12490 471852 12574
rect 472952 12330 473036 12414
rect 520134 12658 520214 12738
rect 520294 12498 520374 12578
rect 520454 12338 520534 12418
rect 475319 12180 475403 12264
rect 520674 12176 520754 12256
rect 476503 12016 476587 12100
rect 478869 11856 478953 11940
rect 480053 11698 480137 11782
rect 520834 12018 520914 12098
rect 520994 11856 521074 11936
rect 521154 11696 521234 11776
rect 482415 11546 482490 11621
rect 521374 11534 521454 11614
rect 483599 11380 483674 11455
rect 485956 11224 486031 11299
rect 487140 11064 487215 11139
rect 521534 11378 521614 11458
rect 521694 11208 521774 11288
rect 521854 11056 521934 11136
rect 489478 10898 489553 10973
rect 522074 10894 522154 10974
rect 490662 10742 490737 10817
rect 493048 10580 493123 10655
rect 494232 10424 494307 10499
rect 522234 10730 522314 10810
rect 522394 10572 522474 10652
rect 522554 10414 522634 10494
rect 496589 10252 496664 10327
rect 522774 10252 522854 10332
rect 497773 10096 497848 10171
rect 500140 9940 500215 10015
rect 501324 9776 501399 9851
rect 522934 10098 523014 10178
rect 523094 9946 523174 10026
rect 523254 9772 523334 9852
rect 503689 9624 503749 9684
rect 523474 9610 523554 9690
rect 504873 9464 504933 9524
rect 507249 9308 507309 9368
rect 508433 9156 508493 9216
rect 523634 9458 523714 9538
rect 549556 373108 552525 376077
rect 563802 260786 563878 260862
rect 524994 256303 525302 256611
rect 563738 256438 563814 256514
rect 563752 254912 563828 254988
rect 524556 253131 524756 253331
rect 524679 252435 525218 252974
rect 562639 244169 563014 244544
rect 558218 170290 558389 170461
rect 523794 9290 523874 9370
rect 523954 9136 524034 9216
rect 510800 8986 510860 9046
rect 524174 8974 524254 9054
rect 511984 8826 512044 8886
rect 514324 8654 514400 8730
rect 515508 8494 515584 8570
rect 524334 8816 524414 8896
rect 524494 8658 524574 8738
rect 524654 8490 524734 8570
rect 517874 8338 517950 8414
rect 524874 8334 524954 8414
rect 519058 8178 519134 8254
rect 521425 8014 521501 8090
rect 522609 7854 522685 7930
rect 525034 8180 525114 8260
rect 548994 151142 549287 151435
rect 549439 150369 549818 150748
rect 558751 73522 558877 73648
rect 525194 8016 525274 8096
rect 539354 7860 539434 7940
rect 524976 7696 525052 7772
rect 539574 7698 539654 7778
rect 526160 7540 526236 7616
rect 528508 7382 528584 7458
rect 529692 7226 529768 7302
rect 539734 7544 539814 7624
rect 539894 7386 539974 7466
rect 540054 7214 540134 7294
rect 532049 7066 532125 7142
rect 540274 7062 540354 7142
rect 533233 6896 533309 6972
rect 535609 6748 535685 6824
rect 536793 6572 536869 6648
rect 540434 6896 540514 6976
rect 550546 54956 550839 55249
rect 540594 6736 540674 6816
rect 550991 54353 551370 54732
rect 540754 6582 540834 6662
rect 539150 6420 539226 6496
rect 565274 6418 565354 6498
rect 540334 6248 540410 6324
rect 542706 6095 542783 6172
rect 543890 5935 543967 6012
rect 565434 6264 565514 6344
rect 565594 6100 565674 6180
rect 565754 5934 565834 6014
rect 546251 5783 546328 5860
rect 566274 5774 566354 5854
rect 547435 5623 547512 5700
rect 549788 5451 549865 5528
rect 550972 5295 551049 5372
rect 566434 5620 566514 5700
rect 566594 5462 566674 5542
rect 566754 5300 566834 5380
rect 553346 5141 553423 5218
rect 567274 5136 567354 5216
rect 554530 4969 554607 5046
rect 556886 4810 556970 4894
rect 558070 4650 558154 4734
rect 567434 4980 567514 5060
rect 567594 4822 567674 4902
rect 567754 4652 567834 4732
rect 560425 4501 560495 4571
rect 568274 4494 568354 4574
rect 561625 4341 561695 4411
rect 563980 4186 564056 4262
rect 565164 4026 565240 4102
rect 568434 4328 568514 4408
rect 568594 4170 568674 4250
rect 577998 353782 580967 356751
rect 568754 4012 568834 4092
rect 567527 3863 567605 3941
rect 569274 3844 569354 3924
rect 568711 3695 568789 3773
rect 569434 3692 569514 3772
rect 569594 3532 569674 3612
rect 569754 3374 569834 3454
rect 570274 3218 570354 3298
rect 570434 3056 570514 3136
rect 570594 2896 570674 2976
rect 570754 2728 570834 2808
rect 571050 3537 571128 3615
rect 572234 3383 572312 3461
rect 574610 3217 574688 3295
rect 575794 3061 575872 3139
rect 578154 2899 578232 2977
rect 579338 2737 579416 2815
<< metal3 >>
rect 16994 703100 21994 705600
rect 68994 703100 73994 705600
rect 120994 703100 125994 705600
rect 166394 703100 171394 705600
rect 171694 703100 173894 704800
rect 174194 703100 176394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 705600
rect 223394 703100 225594 704800
rect 225894 703100 228094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 325094 703100 327294 704800
rect 327594 703100 329794 704800
rect 330094 703100 335094 705600
rect 414194 703100 419194 705600
rect 466194 703100 471194 705600
rect 18574 687352 19364 703100
rect 71019 691045 71393 703100
rect 71019 690671 117078 691045
rect 18574 686562 105509 687352
rect 0 683312 2500 686042
rect 0 682498 101676 683312
rect 0 681042 2500 682498
rect 0 649314 8531 649442
rect 0 644833 3472 649314
rect 8318 644833 8531 649314
rect 0 644642 8531 644833
rect 800 639260 8531 639442
rect 800 634779 3494 639260
rect 8340 634779 8531 639260
rect 800 634642 8531 634779
rect 97764 602175 98028 602176
rect 68712 602055 98030 602175
rect 0 564868 9296 565042
rect 0 560414 4054 564868
rect 9132 560414 9296 564868
rect 0 560242 9296 560414
rect 800 554880 9296 555042
rect 800 550426 4066 554880
rect 9144 550426 9296 554880
rect 800 550242 9296 550426
rect 23187 549740 23547 566272
rect 13230 549380 23547 549740
rect 13230 523750 13590 549380
rect 23667 549032 24027 566262
rect 15964 548672 24027 549032
rect 12603 518260 13733 518566
rect 14039 518260 14045 518566
rect 12772 517330 14156 517650
rect 14476 517330 14482 517650
rect 800 512330 1280 512442
rect 11522 512350 14438 512746
rect 14834 512350 14840 512746
rect 12632 511322 14566 511718
rect 14962 511322 14968 511718
rect 914 511260 1394 511312
rect 0 511174 1394 511260
rect 14388 511174 14652 511180
rect 0 511148 2254 511174
rect 914 511054 2254 511148
rect 1138 510910 2254 511054
rect 12780 510910 14388 511174
rect 14388 510904 14652 510910
rect 800 509966 1280 510078
rect 800 508784 1280 508896
rect 800 507694 1280 507714
rect 800 507602 10048 507694
rect 998 507558 10048 507602
rect 10184 507558 10190 507694
rect 800 506420 2884 506532
rect 2996 506420 9906 506532
rect 10018 506420 10024 506532
rect 15964 480642 16324 548672
rect 17831 511174 18093 511179
rect 17830 511173 26306 511174
rect 17830 510911 17831 511173
rect 18093 510911 26306 511173
rect 17830 510910 26306 510911
rect 17831 510905 18093 510910
rect 13278 480488 16324 480642
rect 13278 480378 16322 480488
rect 12421 475060 24133 475366
rect 24439 475060 24445 475366
rect 12772 474130 24168 474450
rect 24488 474130 24494 474450
rect 0 469108 838 469220
rect 1168 469108 1604 469220
rect 11522 469150 23500 469546
rect 23896 469150 23902 469546
rect 26042 468680 26306 510910
rect 70691 496286 70785 496291
rect 32415 496260 32493 496265
rect 32415 496192 32420 496260
rect 32488 496192 32493 496260
rect 70691 496202 70696 496286
rect 70780 496202 80086 496286
rect 80170 496202 80176 496286
rect 70691 496197 70785 496202
rect 32415 496187 32493 496192
rect 30861 495378 31411 495383
rect 29932 494838 30866 495378
rect 31406 494838 31411 495378
rect 29932 491000 30472 494838
rect 30861 494833 31411 494838
rect 31026 493286 31594 493298
rect 31026 492746 31040 493286
rect 31580 492746 31594 493286
rect 31026 492736 31594 492746
rect 31040 491976 31580 492736
rect 31040 491430 31580 491436
rect 32420 491495 32488 496187
rect 97764 494428 98028 602055
rect 100862 507674 101676 682498
rect 99670 507328 102794 507674
rect 99670 504650 100018 507328
rect 102298 504650 102794 507328
rect 99670 504204 102794 504650
rect 32709 494160 32779 494165
rect 97764 494164 100634 494428
rect 32709 494100 32714 494160
rect 32774 494100 32779 494160
rect 32709 494095 32779 494100
rect 32714 491649 32774 494095
rect 32711 491644 32777 491649
rect 32711 491588 32716 491644
rect 32772 491588 32777 491644
rect 32711 491583 32777 491588
rect 32420 491437 32425 491495
rect 32483 491437 32488 491495
rect 32420 491432 32488 491437
rect 29932 490454 30472 490460
rect 30116 488585 30228 490454
rect 30116 488475 30117 488585
rect 30227 488475 30228 488585
rect 30116 488474 30228 488475
rect 30117 488469 30227 488474
rect 60016 475366 60320 475371
rect 60015 475365 80947 475366
rect 60015 475061 60016 475365
rect 60320 475061 80947 475365
rect 60015 475060 80947 475061
rect 81253 475060 81259 475366
rect 60016 475055 60320 475060
rect 60057 474450 60375 474455
rect 60056 474449 82110 474450
rect 60056 474131 60057 474449
rect 60375 474131 82110 474449
rect 60056 474130 82110 474131
rect 82430 474130 82436 474450
rect 60057 474125 60375 474130
rect 60075 470154 60469 470159
rect 60074 470153 83436 470154
rect 60074 469759 60075 470153
rect 60469 469759 83436 470153
rect 60074 469758 83436 469759
rect 83832 469758 83838 470154
rect 60075 469753 60469 469758
rect 60097 469356 60491 469361
rect 60096 469355 83404 469356
rect 60096 468961 60097 469355
rect 60491 468961 83404 469355
rect 60096 468960 83404 468961
rect 83800 468960 83806 469356
rect 60097 468955 60491 468960
rect 26042 468675 34674 468680
rect 1204 468038 2210 468126
rect 12632 468122 24416 468518
rect 24812 468122 24818 468518
rect 26042 468421 34415 468675
rect 34669 468421 34674 468675
rect 26042 468416 34674 468421
rect 800 467926 2210 468038
rect 1204 467862 2210 467926
rect 1946 467710 2210 467862
rect 12708 467969 33970 467974
rect 12708 467715 33711 467969
rect 33965 467715 33970 467969
rect 12708 467710 33970 467715
rect 800 466744 1280 466856
rect 800 465562 1280 465674
rect 1208 464492 1450 464598
rect 3498 464492 3610 464498
rect 800 464380 3498 464492
rect 1208 464186 1450 464380
rect 3498 464374 3610 464380
rect 800 463198 1988 463310
rect 2100 463198 95464 463310
rect 95576 463198 95582 463310
rect 12730 437437 28906 437442
rect 12730 437183 28647 437437
rect 28901 437183 28906 437437
rect 12730 437178 28906 437183
rect 80599 436423 80905 436429
rect 29695 436117 80599 436423
rect 29695 432166 30001 436117
rect 80599 436111 80905 436117
rect 12615 431860 30001 432166
rect 30350 435514 80692 435834
rect 81012 435514 81018 435834
rect 30350 431250 30670 435514
rect 12768 430930 30670 431250
rect 31070 434810 80686 435206
rect 81082 434810 81088 435206
rect 31070 426346 31466 434810
rect 80710 434560 81106 434566
rect 1061 425998 1444 426125
rect 0 425886 1444 425998
rect 11522 425950 31466 426346
rect 31832 434164 80710 434560
rect 1061 425840 1444 425886
rect 31832 425318 32228 434164
rect 80710 434158 81106 434164
rect 55445 426223 55655 426228
rect 55445 426023 55450 426223
rect 55650 426023 80470 426223
rect 80670 426023 80676 426223
rect 55445 426018 55655 426023
rect 1204 424816 2210 424948
rect 12632 424922 32228 425318
rect 800 424704 2210 424816
rect 55421 424901 55631 424906
rect 1204 424684 2210 424704
rect 1946 424510 2210 424684
rect 12780 424769 32562 424774
rect 12780 424515 32303 424769
rect 32557 424515 32562 424769
rect 55421 424701 55426 424901
rect 55626 424701 80486 424901
rect 80686 424701 80692 424901
rect 55421 424696 55631 424701
rect 12780 424510 32562 424515
rect 55423 424596 55633 424601
rect 55423 424396 55428 424596
rect 55628 424396 80480 424596
rect 80680 424396 80686 424596
rect 55423 424391 55633 424396
rect 800 423522 1280 423634
rect 800 422340 1280 422452
rect 1165 421270 1402 421331
rect 800 421158 2992 421270
rect 3104 421158 3110 421270
rect 1165 421084 1402 421158
rect 5048 420088 5160 420094
rect 800 419976 1780 420088
rect 1892 419976 5048 420088
rect 5048 419970 5160 419976
rect 37903 412914 38113 412919
rect 37903 412714 37908 412914
rect 38108 412714 80418 412914
rect 80618 412714 80624 412914
rect 37903 412709 38113 412714
rect 100370 394242 100634 494164
rect 104719 448630 105509 686562
rect 103912 448182 106444 448630
rect 103912 446394 104310 448182
rect 106146 446394 106444 448182
rect 103912 446048 106444 446394
rect 13278 393978 100634 394242
rect 26147 393365 83873 393671
rect 84179 393365 84185 393671
rect 26147 388966 26453 393365
rect 12767 388660 26453 388966
rect 26992 392834 83834 393154
rect 84154 392834 84160 393154
rect 26992 388050 27312 392834
rect 12714 387730 27312 388050
rect 27916 392236 83820 392632
rect 84216 392236 84222 392632
rect 27916 383146 28312 392236
rect 0 382664 1318 382776
rect 11522 382750 28312 383146
rect 28872 391468 83826 391864
rect 84222 391468 84228 391864
rect 28872 382118 29268 391468
rect 77158 390546 77222 390552
rect 77158 390476 77222 390482
rect 12632 381722 29268 382118
rect 800 381574 1280 381594
rect 800 381482 2222 381574
rect 1270 381310 2222 381482
rect 12780 381569 33392 381574
rect 12780 381315 32967 381569
rect 33221 381315 33392 381569
rect 12780 381310 33392 381315
rect 800 380300 1280 380412
rect 800 379118 1280 379230
rect 0 377936 38866 378048
rect 0 376754 1810 376866
rect 1922 376754 16168 376866
rect 16280 376754 16286 376866
rect 13160 350808 23290 350842
rect 13160 350708 23112 350808
rect 23212 350708 23290 350808
rect 13160 350578 23290 350708
rect 12531 345260 15949 345566
rect 16255 345260 16261 345566
rect 12760 344330 15964 344650
rect 16284 344330 16290 344650
rect 24084 340870 28370 340970
rect 28470 340870 28476 340970
rect 0 339442 1452 339554
rect 11522 339350 15408 339746
rect 15804 339350 15810 339746
rect 800 338362 1280 338372
rect 800 338260 2210 338362
rect 12632 338322 16244 338718
rect 16640 338322 16646 338718
rect 1270 338098 2210 338260
rect 1946 337910 2210 338098
rect 12720 337910 16472 338174
rect 800 337078 1280 337190
rect 800 335896 1280 336008
rect 13964 334826 14076 334832
rect 800 334714 13964 334826
rect 13964 334708 14076 334714
rect 800 333532 2154 333644
rect 2266 333532 14124 333644
rect 14236 333532 14242 333644
rect 13180 307378 15156 307642
rect 15420 307378 15426 307642
rect 12619 302060 13889 302366
rect 14195 302060 14201 302366
rect 12772 301130 14130 301450
rect 14450 301130 14456 301450
rect 0 296220 1430 296332
rect 11522 296150 13166 296546
rect 13562 296150 13568 296546
rect 16208 295878 16472 337910
rect 24084 331439 24184 340870
rect 38766 332004 38866 377936
rect 69415 376866 69525 376871
rect 69414 376865 72878 376866
rect 69414 376755 69415 376865
rect 69525 376755 72878 376865
rect 69414 376754 72878 376755
rect 72990 376754 72996 376866
rect 69415 376749 69525 376754
rect 71906 352176 72018 352182
rect 40082 334978 40598 334983
rect 40082 334472 40087 334978
rect 40593 334472 44239 334978
rect 44745 334472 44751 334978
rect 40082 334467 40598 334472
rect 40074 334060 40566 334065
rect 40074 333578 40079 334060
rect 40561 333578 44253 334060
rect 44735 333578 44741 334060
rect 40074 333573 40566 333578
rect 38761 331999 38871 332004
rect 38761 331899 38766 331999
rect 38866 331899 38871 331999
rect 38761 331894 38871 331899
rect 24327 331439 24437 331444
rect 24084 331339 24332 331439
rect 24432 331339 24437 331439
rect 24327 331334 24437 331339
rect 16765 307642 17027 307647
rect 16764 307641 23326 307642
rect 16764 307379 16765 307641
rect 17027 307520 23326 307641
rect 17027 307420 23124 307520
rect 23224 307420 23326 307520
rect 17027 307379 23326 307420
rect 16764 307378 23326 307379
rect 16765 307373 17027 307378
rect 16208 295823 32738 295878
rect 16208 295645 32495 295823
rect 32673 295645 32738 295823
rect 16208 295614 32738 295645
rect 1172 295150 2210 295152
rect 800 295038 2210 295150
rect 12632 295122 13890 295518
rect 14286 295122 14292 295518
rect 1172 294888 2210 295038
rect 1946 294710 2210 294888
rect 12780 294917 32094 294974
rect 12780 294739 31883 294917
rect 32061 294739 32094 294917
rect 12780 294710 32094 294739
rect 800 293856 1280 293968
rect 800 292674 1280 292786
rect 71906 291604 72018 352064
rect 800 291492 72018 291604
rect 800 290310 2144 290422
rect 2256 290310 5902 290422
rect 5748 281740 5860 290310
rect 40648 285265 42248 285270
rect 40648 283675 40653 285265
rect 42243 283675 66377 285265
rect 67967 283675 67973 285265
rect 40648 283670 42248 283675
rect 14880 281877 15184 281882
rect 14879 281876 66223 281877
rect 14879 281740 14880 281876
rect 5748 281628 14880 281740
rect 14879 281572 14880 281628
rect 15184 281572 66223 281876
rect 14879 281571 66223 281572
rect 66529 281571 66535 281877
rect 14880 281566 15184 281571
rect 15609 281134 15938 281138
rect 15609 281133 66290 281134
rect 15609 280815 15615 281133
rect 15933 280815 66290 281133
rect 15614 280814 66290 280815
rect 66610 280814 66616 281134
rect 77160 279536 77220 390476
rect 77941 389988 78075 389993
rect 77940 389987 78076 389988
rect 77940 389853 77941 389987
rect 78075 389853 78076 389987
rect 77158 279530 77222 279536
rect 77158 279460 77222 279466
rect 77940 279088 78076 389853
rect 78789 389350 79199 389355
rect 14274 278824 78076 279088
rect 78788 389349 79200 389350
rect 78788 388939 78789 389349
rect 79199 388939 79200 389349
rect 14274 264642 14538 278824
rect 77152 278282 77158 278346
rect 77222 278282 77228 278346
rect 45652 277951 47252 277956
rect 45652 276361 45657 277951
rect 47247 276361 66317 277951
rect 67907 276361 67913 277951
rect 45652 276356 47252 276361
rect 12824 264378 14538 264642
rect 12755 259060 14879 259366
rect 15185 259060 15191 259366
rect 12614 258130 15614 258450
rect 15934 258130 15940 258450
rect 1102 253310 1512 253320
rect 0 253198 1512 253310
rect 1102 253188 1512 253198
rect 11522 253150 15582 253546
rect 15978 253150 15984 253546
rect 1270 252128 2210 252138
rect 800 252016 2210 252128
rect 12632 252122 14736 252518
rect 15132 252122 15138 252518
rect 1270 251874 2210 252016
rect 1946 251710 2210 251874
rect 12780 251710 14090 251974
rect 800 250834 1280 250946
rect 800 249652 1280 249764
rect 800 248470 12314 248582
rect 11476 247400 11588 247406
rect 800 247288 2464 247400
rect 2576 247288 11476 247400
rect 11476 247282 11588 247288
rect 0 220396 9632 220488
rect 0 215890 4310 220396
rect 9440 215890 9632 220396
rect 12202 220120 12314 248470
rect 13880 248558 14080 251710
rect 13880 248358 25064 248558
rect 13573 247400 13683 247405
rect 13572 247399 23502 247400
rect 13572 247289 13573 247399
rect 13683 247289 23502 247399
rect 13572 247288 23502 247289
rect 13573 247283 13683 247288
rect 23390 224272 23502 247288
rect 23390 224160 24984 224272
rect 24872 223860 24984 224160
rect 61926 224204 62598 224209
rect 61926 223860 61931 224204
rect 24872 223748 61931 223860
rect 61926 223542 61931 223748
rect 62593 223542 69747 224204
rect 70409 223542 70415 224204
rect 61926 223537 62598 223542
rect 45942 223392 46614 223397
rect 39307 223387 45947 223392
rect 39307 222735 39312 223387
rect 39964 222735 45947 223387
rect 39307 222730 45947 222735
rect 46609 222730 46614 223392
rect 45942 222725 46614 222730
rect 61872 223392 62544 223397
rect 61872 222730 61877 223392
rect 62539 222730 69873 223392
rect 70535 222730 70541 223392
rect 61872 222725 62544 222730
rect 77160 220120 77220 278282
rect 12202 220008 77220 220120
rect 0 215688 9632 215890
rect 800 210358 9632 210488
rect 800 205852 4284 210358
rect 9414 205852 9632 210358
rect 800 205688 9632 205852
rect 0 178310 9505 178488
rect 0 173829 3756 178310
rect 8602 173829 9505 178310
rect 0 173688 9505 173829
rect 800 168320 9505 168488
rect 800 163839 3676 168320
rect 8522 163839 9505 168320
rect 800 163688 9505 163839
rect 78788 137220 79200 388939
rect 79990 388351 80235 388356
rect 13614 136960 79200 137220
rect 79989 388350 80236 388351
rect 79989 388105 79990 388350
rect 80235 388105 80236 388350
rect 13614 136956 79080 136960
rect 44018 133617 45139 133622
rect 44018 132506 44023 133617
rect 45134 132506 78004 133617
rect 79115 132506 79121 133617
rect 44018 132501 45139 132506
rect 13381 131638 22349 131944
rect 22655 131638 22661 131944
rect 50118 131546 50506 131551
rect 50118 131168 50123 131546
rect 50501 131168 78265 131546
rect 78643 131168 78649 131546
rect 50118 131163 50506 131168
rect 23322 131028 23642 131034
rect 13336 130708 23322 131028
rect 23322 130702 23642 130708
rect 42538 130801 42650 130806
rect 42538 130699 42543 130801
rect 42645 130699 42650 130801
rect 994 125688 1590 125821
rect 12086 125728 23176 126124
rect 23572 125728 23578 126124
rect 0 125576 1590 125688
rect 994 125450 1590 125576
rect 13196 124700 23194 125096
rect 23590 124700 23596 125096
rect 1270 124506 2774 124552
rect 800 124394 2774 124506
rect 1270 124288 2774 124394
rect 800 123212 1280 123324
rect 42538 122414 42650 130699
rect 50092 129165 50480 129170
rect 50092 128787 50097 129165
rect 50475 128787 78253 129165
rect 78631 128787 78637 129165
rect 50092 128782 50480 128787
rect 44567 127856 45688 127861
rect 44567 126745 44572 127856
rect 45683 126745 47794 127856
rect 48905 126745 48911 127856
rect 44567 126740 45688 126745
rect 11188 122302 42650 122414
rect 800 122030 1280 122142
rect 11188 120960 11300 122302
rect 800 120848 11300 120960
rect 800 119666 1558 119778
rect 1678 119666 77898 119778
rect 78010 119666 78016 119778
rect 79989 94116 80236 388105
rect 116704 347944 117078 690671
rect 115878 347766 118262 347944
rect 115878 345626 116072 347766
rect 118072 345626 118262 347766
rect 115878 345460 118262 345626
rect 122792 287156 123728 703100
rect 168369 697685 168783 703100
rect 146740 697271 168783 697685
rect 128832 655062 132832 658652
rect 128832 653816 130007 655062
rect 131253 653816 132832 655062
rect 128832 614289 132832 653816
rect 128832 612731 130013 614289
rect 131571 612731 132832 614289
rect 126591 591465 127549 596408
rect 128832 595370 132832 612731
rect 136832 657462 140832 658478
rect 136832 656216 138173 657462
rect 139419 656216 140832 657462
rect 136832 644370 140832 656216
rect 136832 639691 136986 644370
rect 140674 639691 140832 644370
rect 136832 598903 140832 639691
rect 136832 597505 137993 598903
rect 139391 597505 140832 598903
rect 126591 591344 126893 591465
rect 127014 591344 127549 591465
rect 126591 496285 127549 591344
rect 128823 595069 132844 595370
rect 128823 589599 129074 595069
rect 132598 589599 132844 595069
rect 128823 589258 132844 589599
rect 126591 496203 127105 496285
rect 127187 496203 127549 496285
rect 121856 286830 124852 287156
rect 121856 284192 122182 286830
rect 124562 284192 124852 286830
rect 121856 283880 124852 284192
rect 126591 276719 127549 496203
rect 13645 93869 80236 94116
rect 124735 275761 127549 276719
rect 128832 565062 132832 589258
rect 128832 563816 130007 565062
rect 131253 564299 132832 565062
rect 128832 563101 130223 563816
rect 131421 563101 132832 564299
rect 128832 520558 132832 563101
rect 128832 520254 130494 520558
rect 130798 520254 132832 520558
rect 128832 490999 132832 520254
rect 128832 490461 130371 490999
rect 130909 490461 132832 490999
rect 128832 481602 132832 490461
rect 128832 481298 130662 481602
rect 130966 481298 132832 481602
rect 128832 478334 132832 481298
rect 128832 472030 129018 478334
rect 132644 472030 132832 478334
rect 128832 463309 132832 472030
rect 128832 463199 130729 463309
rect 130839 463199 132832 463309
rect 128832 436422 132832 463199
rect 128832 436118 130708 436422
rect 131012 436118 132832 436422
rect 128832 424595 132832 436118
rect 128832 424397 130461 424595
rect 130659 424397 132832 424595
rect 128832 412913 132832 424397
rect 128832 412715 130591 412913
rect 130789 412715 132832 412913
rect 128832 393670 132832 412715
rect 128832 393366 130804 393670
rect 131108 393366 132832 393670
rect 128832 385062 132832 393366
rect 128832 383816 130159 385062
rect 131405 383816 132832 385062
rect 128832 380144 132832 383816
rect 128832 379827 128918 380144
rect 132762 379827 132832 380144
rect 128832 377026 132832 379827
rect 128832 376582 128962 377026
rect 132722 376582 132832 377026
rect 128832 364692 132832 376582
rect 128832 363838 128893 364692
rect 132628 363838 132832 364692
rect 128832 356126 132832 363838
rect 128832 355822 130472 356126
rect 130776 355822 132832 356126
rect 128832 334977 132832 355822
rect 128832 334473 130656 334977
rect 131160 334473 132832 334977
rect 128832 310649 132832 334473
rect 128832 310102 128934 310649
rect 132738 310102 132832 310649
rect 128832 302365 132832 310102
rect 128832 302061 130624 302365
rect 130928 302061 132832 302365
rect 128832 295062 132832 302061
rect 128832 293816 129929 295062
rect 131175 293816 132832 295062
rect 128832 279558 132832 293816
rect 128832 279254 130802 279558
rect 131106 279254 132832 279558
rect 13355 88438 29441 88744
rect 29747 88438 29753 88744
rect 29646 87828 29966 87834
rect 13336 87508 29646 87828
rect 29646 87502 29966 87508
rect 984 82466 1294 82602
rect 12086 82528 29596 82924
rect 29992 82528 29998 82924
rect 0 82354 1294 82466
rect 984 82231 1294 82354
rect 29604 81896 30000 81902
rect 13156 81500 29604 81896
rect 29604 81494 30000 81500
rect 1238 81284 2876 81352
rect 800 81172 2876 81284
rect 1238 81088 2876 81172
rect 13220 81088 27430 81352
rect 800 79990 1280 80102
rect 800 78808 1280 78920
rect 800 77626 1280 77738
rect 800 76444 1280 76556
rect 27166 66708 27430 81088
rect 120566 81344 120962 81350
rect 27166 66464 31310 66708
rect 42786 59528 44174 59533
rect 41183 59527 44175 59528
rect 41183 59523 42786 59527
rect 41183 58143 41188 59523
rect 42568 58143 42786 59523
rect 41183 58139 42786 58143
rect 44174 58139 44175 59527
rect 41183 58138 44175 58139
rect 42786 58133 44174 58138
rect 40006 57258 42564 57263
rect 40006 57188 42439 57258
rect 42509 57188 42564 57258
rect 40006 57183 42564 57188
rect 40012 57078 42868 57083
rect 40012 57008 42745 57078
rect 42815 57008 42868 57078
rect 40012 57003 42868 57008
rect 27034 50852 31338 51096
rect 13381 45238 24125 45544
rect 24431 45238 24437 45544
rect 13336 44308 24086 44628
rect 24406 44308 24412 44628
rect 12086 39328 23432 39724
rect 23828 39328 23834 39724
rect 0 39132 1350 39244
rect 13196 38300 23402 38696
rect 23798 38300 23804 38696
rect 27034 38152 27298 50852
rect 120566 41327 120962 80948
rect 120566 40933 120567 41327
rect 120961 40933 120962 41327
rect 120566 40932 120962 40933
rect 120567 40927 120961 40932
rect 1168 38062 2774 38152
rect 800 37950 2774 38062
rect 1168 37888 2774 37950
rect 13340 37888 27298 38152
rect 800 36768 1280 36880
rect 800 35586 1280 35698
rect 1092 34516 1362 34609
rect 0 34404 1362 34516
rect 1092 34319 1362 34404
rect 1131 33334 1362 33416
rect 0 33222 1362 33334
rect 1131 33126 1362 33222
rect 124735 18189 125693 275761
rect 128832 234956 132832 279254
rect 128832 234296 130162 234956
rect 130822 234296 132832 234956
rect 128832 205062 132832 234296
rect 128832 203816 130159 205062
rect 131405 203816 132832 205062
rect 128832 173511 132832 203816
rect 128832 168834 129023 173511
rect 132621 168834 132832 173511
rect 128832 136828 132832 168834
rect 128832 136524 130688 136828
rect 130992 136524 132832 136828
rect 128832 131545 132832 136524
rect 128832 131169 130506 131545
rect 130882 131169 132832 131545
rect 128832 119777 132832 131169
rect 128832 119667 130809 119777
rect 130919 119667 132832 119777
rect 128832 119218 132832 119667
rect 128832 112664 129090 119218
rect 132624 112664 132832 119218
rect 128832 88743 132832 112664
rect 128832 88439 130670 88743
rect 130974 88439 132832 88743
rect 128832 46645 132832 88439
rect 128832 45059 130143 46645
rect 131729 45059 132832 46645
rect 128832 44076 132832 45059
rect 128832 43772 130662 44076
rect 130966 43772 132832 44076
rect 128832 34732 132832 43772
rect 136832 573356 140832 597505
rect 136832 572158 138121 573356
rect 139319 572158 140832 573356
rect 136832 567462 140832 572158
rect 136832 566216 138287 567462
rect 139533 566216 140832 567462
rect 136832 519505 140832 566216
rect 136832 519187 138459 519505
rect 138777 519187 140832 519505
rect 136832 491975 140832 519187
rect 136832 491437 138631 491975
rect 139169 491437 140832 491975
rect 136832 480499 140832 491437
rect 136832 480181 138317 480499
rect 138635 480181 140832 480499
rect 136832 477462 140832 480181
rect 136832 476216 138401 477462
rect 139647 476216 140832 477462
rect 136832 435833 140832 476216
rect 136832 435515 138711 435833
rect 139029 435515 140832 435833
rect 136832 424900 140832 435515
rect 136832 424702 138589 424900
rect 138787 424702 140832 424900
rect 136832 404667 140832 424702
rect 136832 404349 138495 404667
rect 138813 404349 140832 404667
rect 136832 401010 140832 404349
rect 136832 391475 137099 401010
rect 140611 391475 140832 401010
rect 136832 387462 140832 391475
rect 136832 386216 138267 387462
rect 139513 386216 140832 387462
rect 136832 379269 140832 386216
rect 136832 378850 136999 379269
rect 140729 378850 140832 379269
rect 136832 362468 140832 378850
rect 136832 361328 136912 362468
rect 140668 361328 140832 362468
rect 136832 354993 140832 361328
rect 136832 354675 138801 354993
rect 139119 354675 140832 354993
rect 136832 334059 140832 354675
rect 136832 333579 138718 334059
rect 139198 333579 140832 334059
rect 136832 309624 140832 333579
rect 136832 309106 136918 309624
rect 140746 309106 140832 309624
rect 136832 301449 140832 309106
rect 136832 301131 138483 301449
rect 138801 301131 140832 301449
rect 136832 297462 140832 301131
rect 136832 296216 138115 297462
rect 139361 296216 140832 297462
rect 136832 278551 140832 296216
rect 136832 278233 138369 278551
rect 138687 278233 140832 278551
rect 136832 233696 140832 278233
rect 136832 233036 138658 233696
rect 139318 233036 140832 233696
rect 136832 207462 140832 233036
rect 136832 206216 138191 207462
rect 139437 206216 140832 207462
rect 136832 136033 140832 206216
rect 146740 146616 147154 697271
rect 220111 693525 220373 703100
rect 160762 693263 220373 693525
rect 145758 146268 148578 146616
rect 145758 143960 146008 146268
rect 148318 143960 148578 146268
rect 145758 143656 148578 143960
rect 136832 135715 138813 136033
rect 139131 135715 140832 136033
rect 136832 129164 140832 135715
rect 136832 128788 138734 129164
rect 139110 128788 140832 129164
rect 136832 117462 140832 128788
rect 136832 116216 138173 117462
rect 139419 116216 140832 117462
rect 136832 87827 140832 116216
rect 136832 87509 138953 87827
rect 139271 87509 140832 87827
rect 136832 59527 140832 87509
rect 160762 66334 161024 693263
rect 331404 680832 331796 703100
rect 415856 686754 416308 703100
rect 467586 686834 468038 703100
rect 511394 698944 516194 705600
rect 511394 693868 511510 698944
rect 516020 693868 516194 698944
rect 511394 693672 516194 693868
rect 521394 698932 526194 705600
rect 567394 703100 572394 705600
rect 521394 693856 521554 698932
rect 526064 693856 526194 698932
rect 521394 693672 526194 693856
rect 415856 686302 427878 686754
rect 331404 680440 424246 680832
rect 423854 607278 424246 680440
rect 422464 606998 426030 607278
rect 422464 604042 422844 606998
rect 425668 604042 426030 606998
rect 422464 603712 426030 604042
rect 427426 430644 427878 686302
rect 430574 686382 468038 686834
rect 426340 430286 428862 430644
rect 426340 428204 426592 430286
rect 428498 428204 428862 430286
rect 426340 427878 428862 428204
rect 427838 287992 428290 287995
rect 430574 287992 431026 686382
rect 467586 686276 468038 686382
rect 568648 683460 569100 703100
rect 433826 683008 569100 683460
rect 426826 287604 431158 287992
rect 426826 284006 427136 287604
rect 430734 284006 431158 287604
rect 426826 283660 431158 284006
rect 433826 200154 434278 683008
rect 583100 680372 585600 683784
rect 436838 679920 585600 680372
rect 436838 200154 437290 679920
rect 583100 678784 585600 679920
rect 444177 657462 448177 658360
rect 444177 656216 445405 657462
rect 446651 656216 448177 657462
rect 444177 640383 448177 656216
rect 444177 635697 444374 640383
rect 448011 635697 448177 640383
rect 444177 599100 448177 635697
rect 444177 598724 445990 599100
rect 446366 598724 448177 599100
rect 444177 592191 448177 598724
rect 444177 591873 445999 592191
rect 446317 591873 448177 592191
rect 444177 567462 448177 591873
rect 444177 566216 445481 567462
rect 446727 566216 448177 567462
rect 444177 516489 448177 566216
rect 444177 516171 446115 516489
rect 446433 516171 448177 516489
rect 444177 511391 448177 516171
rect 444177 511073 445899 511391
rect 446217 511073 448177 511391
rect 444177 495191 448177 511073
rect 444177 494873 445837 495191
rect 446155 494873 448177 495191
rect 444177 492461 448177 494873
rect 444177 492239 445803 492461
rect 446025 492239 448177 492461
rect 444177 482287 448177 492239
rect 444177 481969 445789 482287
rect 446107 481969 448177 482287
rect 444177 477462 448177 481969
rect 444177 476216 445367 477462
rect 446613 476216 448177 477462
rect 444177 387462 448177 476216
rect 452177 655062 456177 658558
rect 452177 653816 453593 655062
rect 454839 653816 456177 655062
rect 452177 598226 456177 653816
rect 573658 645170 584800 645384
rect 573658 640732 573828 645170
rect 578952 640732 584800 645170
rect 573658 640584 584800 640732
rect 573658 635200 585600 635384
rect 573658 630762 573842 635200
rect 578966 630762 585600 635200
rect 573658 630584 585600 630762
rect 538246 615607 540250 615612
rect 493997 613613 538251 615607
rect 540245 613613 540250 615607
rect 493997 606979 495991 613613
rect 538246 613608 540250 613613
rect 583264 611666 583348 611671
rect 583264 611592 583269 611666
rect 583343 611592 583348 611666
rect 583264 611587 583348 611592
rect 541054 608974 543058 608979
rect 493997 604979 495991 604985
rect 498783 606980 541059 608974
rect 543053 606980 543058 608974
rect 452177 597850 453800 598226
rect 454176 597850 456177 598226
rect 452177 593107 456177 597850
rect 498783 597333 500777 606980
rect 541054 606975 543058 606980
rect 560286 603833 560674 603838
rect 509743 603455 509749 603833
rect 510127 603455 560291 603833
rect 560669 603455 560674 603833
rect 560286 603450 560674 603455
rect 561258 602873 561646 602878
rect 509791 602495 509797 602873
rect 510175 602495 561263 602873
rect 561641 602495 561646 602873
rect 561258 602490 561646 602495
rect 540022 598379 571260 598384
rect 540022 598125 540027 598379
rect 540281 598125 571260 598379
rect 540022 598120 571260 598125
rect 498783 595333 500777 595339
rect 452177 592803 454030 593107
rect 454334 592803 456177 593107
rect 452177 565062 456177 592803
rect 564583 592802 564589 593108
rect 564895 592802 571819 593108
rect 564644 591872 564650 592192
rect 564970 591872 571832 592192
rect 583269 589199 583343 611587
rect 584048 599628 584160 599634
rect 584048 590684 584160 599516
rect 584048 590384 584160 590572
rect 584048 590272 585600 590384
rect 584048 589199 585600 589202
rect 583269 589125 585600 589199
rect 584048 589090 585600 589125
rect 584320 587908 584800 588020
rect 564504 586892 564510 587288
rect 564906 586892 573030 587288
rect 584320 586726 584800 586838
rect 564422 585864 564428 586260
rect 564824 585864 571886 586260
rect 582258 585656 584408 585716
rect 563360 585567 563456 585572
rect 563360 585481 563365 585567
rect 563451 585481 571745 585567
rect 582258 585544 584800 585656
rect 563360 585476 563456 585481
rect 582258 585452 584408 585544
rect 584286 584362 585600 584474
rect 452177 563816 453515 565062
rect 454761 563816 456177 565062
rect 452177 515597 456177 563816
rect 575498 556038 584800 556162
rect 575498 551600 575644 556038
rect 580768 551600 584800 556038
rect 575498 551362 584800 551600
rect 575498 546004 585600 546162
rect 575498 541566 575630 546004
rect 580754 541566 585600 546004
rect 575498 541362 585600 541566
rect 523947 528823 523953 529377
rect 524507 528823 536228 529377
rect 524032 528018 524038 528338
rect 524358 528018 535555 528338
rect 524160 527410 524166 527730
rect 524486 527410 535105 527730
rect 534105 526846 534666 526880
rect 524144 526285 524150 526846
rect 524711 526285 534666 526846
rect 534105 524792 534666 526285
rect 534785 524792 535105 527410
rect 535235 524792 535555 528018
rect 535674 524792 536228 528823
rect 452177 515279 454037 515597
rect 454355 515279 456177 515597
rect 452177 512307 456177 515279
rect 551778 517320 571440 517584
rect 551778 512602 552042 517320
rect 540072 512597 552042 512602
rect 540072 512343 540077 512597
rect 540331 512343 552042 512597
rect 540072 512338 552042 512343
rect 452177 512003 453982 512307
rect 454286 512003 456177 512307
rect 452177 496107 456177 512003
rect 561361 512002 561367 512308
rect 561673 512002 571813 512308
rect 561430 511072 561436 511392
rect 561756 511072 571922 511392
rect 561328 506092 561334 506488
rect 561730 506092 572996 506488
rect 561376 505064 561382 505460
rect 561778 505064 571930 505460
rect 574832 503932 574992 504772
rect 582266 504652 583162 504916
rect 583426 504652 583432 504916
rect 574832 503772 582282 503932
rect 582442 503772 582448 503932
rect 559842 502678 559848 502790
rect 559960 502678 582848 502790
rect 452177 495803 453846 496107
rect 454150 495803 456177 496107
rect 452177 490003 456177 495803
rect 452177 489805 454027 490003
rect 454225 489805 456177 490003
rect 452177 483340 456177 489805
rect 452177 483036 454076 483340
rect 454380 483036 456177 483340
rect 452177 475062 456177 483036
rect 452177 473816 453439 475062
rect 454685 473816 456177 475062
rect 451716 390552 451776 390602
rect 451714 390546 451778 390552
rect 451714 390476 451778 390482
rect 451236 389988 451372 389994
rect 450424 389350 450836 389356
rect 442634 387140 443287 387242
rect 442628 386487 442634 387140
rect 443287 386487 443293 387140
rect 439833 385423 439963 385526
rect 439337 383259 439555 383426
rect 438563 382473 438742 382692
rect 438563 381382 438742 382294
rect 439337 381480 439555 383041
rect 439332 381475 439560 381480
rect 438558 381377 438747 381382
rect 438558 381198 438563 381377
rect 438742 381198 438747 381377
rect 439332 381257 439337 381475
rect 439555 381257 439560 381475
rect 439833 381390 439963 385293
rect 441444 384588 442145 384776
rect 441444 381757 442145 383887
rect 441439 381752 442150 381757
rect 439332 381252 439560 381257
rect 439828 381385 439968 381390
rect 439828 381255 439833 381385
rect 439963 381255 439968 381385
rect 439828 381250 439968 381255
rect 438558 381193 438747 381198
rect 441439 381051 441444 381752
rect 442145 381051 442150 381752
rect 442634 381677 443287 386487
rect 444177 386216 445481 387462
rect 446727 386216 448177 387462
rect 441439 381046 442150 381051
rect 442629 381672 443292 381677
rect 442629 381019 442634 381672
rect 443287 381019 443292 381672
rect 442629 381014 443292 381019
rect 444177 317191 448177 386216
rect 449325 388351 449759 388357
rect 449325 375122 449759 387917
rect 450424 376426 450836 388938
rect 451236 381275 451372 389852
rect 451716 382218 451776 390476
rect 452177 385062 456177 473816
rect 452177 383816 453515 385062
rect 454761 383816 456177 385062
rect 451711 382213 451781 382218
rect 451711 382153 451716 382213
rect 451776 382153 451781 382213
rect 451711 382148 451781 382153
rect 451231 381270 451377 381275
rect 451231 381134 451236 381270
rect 451372 381134 451377 381270
rect 451231 381129 451377 381134
rect 450419 376421 450841 376426
rect 450419 376009 450424 376421
rect 450836 376009 450841 376421
rect 450419 376004 450841 376009
rect 452177 376076 456177 383816
rect 461190 502082 581544 502194
rect 461190 377385 461302 502082
rect 533948 501689 534044 501694
rect 533948 501603 533953 501689
rect 534039 501684 563451 501689
rect 534039 501608 563370 501684
rect 563446 501608 563451 501684
rect 534039 501603 563451 501608
rect 533948 501598 534044 501603
rect 533960 501247 534056 501252
rect 533960 501161 533965 501247
rect 534051 501161 571303 501247
rect 533960 501156 534056 501161
rect 581432 499780 581544 502082
rect 582736 500962 582848 502678
rect 582736 500850 584088 500962
rect 584200 500850 585600 500962
rect 584288 499780 584508 499829
rect 581432 499668 585600 499780
rect 584288 499598 584508 499668
rect 584320 498486 584800 498598
rect 584320 497304 584800 497416
rect 583162 496279 584404 496280
rect 561165 495802 561171 496108
rect 561477 495802 571855 496108
rect 583157 496017 583163 496279
rect 583425 496234 584404 496279
rect 583425 496122 584800 496234
rect 583425 496017 584404 496122
rect 583162 496016 584404 496017
rect 561234 494872 561240 495192
rect 561560 494872 571746 495192
rect 584270 494940 585600 495052
rect 543806 492462 544030 492468
rect 542206 490004 542406 490010
rect 528276 488997 528282 489426
rect 528711 488997 533179 489426
rect 542206 488836 542406 489804
rect 542201 488831 542411 488836
rect 542201 488631 542206 488831
rect 542406 488631 542411 488831
rect 542201 488626 542411 488631
rect 543806 484869 544030 492238
rect 560784 489892 560790 490288
rect 561186 489892 572996 490288
rect 560716 488864 560722 489260
rect 561118 488864 571886 489260
rect 561774 488716 561780 488776
rect 561746 488452 561780 488716
rect 561774 488448 561780 488452
rect 562108 488716 562114 488776
rect 562108 488452 571864 488716
rect 582308 488452 583194 488716
rect 583458 488452 583464 488716
rect 562108 488448 562114 488452
rect 550026 488260 550122 488265
rect 550026 488174 550031 488260
rect 550117 488174 558691 488260
rect 550026 488169 550122 488174
rect 558605 485997 558691 488174
rect 581531 485997 581617 486003
rect 558605 485911 581531 485997
rect 581531 485905 581617 485911
rect 541480 484645 544030 484869
rect 570050 484520 571364 484784
rect 487304 480710 487700 480716
rect 486350 479452 486746 479458
rect 486350 472659 486746 479056
rect 487304 473687 487700 480314
rect 537940 477407 538369 481287
rect 562984 479508 563288 479513
rect 556413 479202 556419 479508
rect 556725 479507 563289 479508
rect 556725 479203 562984 479507
rect 563288 479203 563289 479507
rect 556725 479202 563289 479203
rect 562984 479197 563288 479202
rect 563127 478592 563445 478597
rect 556608 478272 556614 478592
rect 556934 478591 563446 478592
rect 556934 478273 563127 478591
rect 563445 478273 563446 478591
rect 556934 478272 563446 478273
rect 563127 478267 563445 478272
rect 537940 476972 538369 476978
rect 487304 473293 487305 473687
rect 487699 473293 487700 473687
rect 487304 473292 487700 473293
rect 487305 473287 487699 473292
rect 486350 472265 486351 472659
rect 486745 472265 486746 472659
rect 486350 472264 486746 472265
rect 486351 472259 486745 472264
rect 483617 471076 483727 471081
rect 461910 471075 483728 471076
rect 461910 470965 483617 471075
rect 483727 470965 483728 471075
rect 461910 470964 483728 470965
rect 461910 377751 462022 470964
rect 483617 470959 483727 470964
rect 570052 470762 570289 484520
rect 570853 479202 570859 479508
rect 571165 479380 571721 479508
rect 571165 479379 583864 479380
rect 571165 479269 583753 479379
rect 583863 479269 583869 479379
rect 571165 479268 583864 479269
rect 571165 479202 571721 479268
rect 570846 478272 570852 478592
rect 571172 478272 572030 478592
rect 570698 473292 570704 473688
rect 571100 473292 572996 473688
rect 570714 472264 570720 472660
rect 571116 472264 571894 472660
rect 576384 471330 576621 472116
rect 581956 471852 582282 472116
rect 582546 471852 582552 472116
rect 576384 471093 579494 471330
rect 570052 470525 578798 470762
rect 461910 377649 461915 377751
rect 462017 377649 462022 377751
rect 461910 377644 462022 377649
rect 505921 390521 506251 390527
rect 461190 377283 461195 377385
rect 461297 377283 461302 377385
rect 461190 377278 461302 377283
rect 505921 377156 506251 390191
rect 517539 388631 517685 388636
rect 517539 388495 517544 388631
rect 517680 388626 520548 388631
rect 517680 388500 520417 388626
rect 520543 388500 520548 388626
rect 517680 388495 520548 388500
rect 517539 388490 517685 388495
rect 517551 387928 517697 387933
rect 517551 387792 517556 387928
rect 517692 387923 520270 387928
rect 517692 387797 520139 387923
rect 520265 387797 520270 387923
rect 517692 387792 520270 387797
rect 517551 387787 517697 387792
rect 517683 386264 517829 386269
rect 517683 386128 517688 386264
rect 517824 386259 519240 386264
rect 517824 386133 519109 386259
rect 519235 386133 519240 386259
rect 517824 386128 519240 386133
rect 517683 386123 517829 386128
rect 517521 385247 517667 385252
rect 517521 385111 517526 385247
rect 517662 385242 520222 385247
rect 517662 385116 520091 385242
rect 520217 385116 520222 385242
rect 517662 385111 520222 385116
rect 517521 385106 517667 385111
rect 578561 383388 578798 470525
rect 516800 383269 516884 383274
rect 516800 383195 516805 383269
rect 516879 383264 520865 383269
rect 516879 383200 520796 383264
rect 520860 383200 520865 383264
rect 516879 383195 520865 383200
rect 516800 383190 516884 383195
rect 564181 383151 578798 383388
rect 506917 380963 506987 380968
rect 521195 380963 521261 380966
rect 506917 380903 506922 380963
rect 506982 380961 521261 380963
rect 506982 380905 521200 380961
rect 521256 380905 521261 380961
rect 506982 380903 521261 380905
rect 506917 380898 506987 380903
rect 521195 380900 521261 380903
rect 516865 378844 516935 378849
rect 519141 378844 519207 378847
rect 516865 378784 516870 378844
rect 516930 378842 519207 378844
rect 516930 378786 519146 378842
rect 519202 378786 519207 378842
rect 516930 378784 519207 378786
rect 516865 378779 516935 378784
rect 519141 378781 519207 378784
rect 516816 378596 516920 378601
rect 516816 378502 516821 378596
rect 516915 378591 519179 378596
rect 516915 378507 519090 378591
rect 519174 378507 519179 378591
rect 516915 378502 519179 378507
rect 516816 378497 516920 378502
rect 516876 378368 516980 378373
rect 516876 378274 516881 378368
rect 516975 378363 519239 378368
rect 516975 378279 519150 378363
rect 519234 378279 519239 378363
rect 516975 378274 519239 378279
rect 516876 378269 516980 378274
rect 516948 378086 517052 378091
rect 516948 377992 516953 378086
rect 517047 378081 519379 378086
rect 517047 377997 519290 378081
rect 519374 377997 519379 378081
rect 517047 377992 519379 377997
rect 516948 377987 517052 377992
rect 505916 377151 506256 377156
rect 505916 376821 505921 377151
rect 506251 376821 506256 377151
rect 505916 376816 506256 376821
rect 549551 376077 552530 376082
rect 449312 375111 449774 375122
rect 449312 374677 449325 375111
rect 449759 374677 449774 375111
rect 449312 374668 449774 374677
rect 444177 316873 446017 317191
rect 446335 316873 448177 317191
rect 444177 310980 448177 316873
rect 444177 301612 444618 310980
rect 447812 301612 448177 310980
rect 444177 297680 448177 301612
rect 444174 297462 448177 297680
rect 444174 296624 445367 297462
rect 444177 296216 445367 296624
rect 446613 296216 448177 297462
rect 444177 277991 448177 296216
rect 444177 277673 446021 277991
rect 446339 277673 448177 277991
rect 444177 244543 448177 277673
rect 444177 244170 445726 244543
rect 446099 244170 448177 244543
rect 444177 207462 448177 244170
rect 444177 206216 445597 207462
rect 446843 206216 448177 207462
rect 433855 167330 434271 200154
rect 431050 167041 434772 167330
rect 431050 163637 431353 167041
rect 434495 163637 434772 167041
rect 431050 163361 434772 163637
rect 436856 68598 437272 200154
rect 444177 180774 448177 206216
rect 444177 179958 444303 180774
rect 448071 179958 448177 180774
rect 444177 117462 448177 179958
rect 452177 373109 452461 376076
rect 455428 373109 456177 376076
rect 452177 318107 456177 373109
rect 545324 373108 545330 376077
rect 548299 373108 549556 376077
rect 552525 373108 552530 376077
rect 549551 373103 552530 373108
rect 490953 349378 491099 349383
rect 490953 349242 490958 349378
rect 491094 349350 521286 349378
rect 491094 349270 521154 349350
rect 521234 349270 521286 349350
rect 491094 349242 521286 349270
rect 490953 349237 491099 349242
rect 490901 349058 491047 349063
rect 490901 348922 490906 349058
rect 491042 349040 521104 349058
rect 491042 348960 520994 349040
rect 521074 348960 521104 349040
rect 491042 348922 521104 348960
rect 490901 348917 491047 348922
rect 490885 348720 491031 348725
rect 490885 348584 490890 348720
rect 491026 348700 520934 348720
rect 491026 348620 520834 348700
rect 520914 348620 520934 348700
rect 491026 348584 520934 348620
rect 490885 348579 491031 348584
rect 490953 348366 491099 348371
rect 490953 348230 490958 348366
rect 491094 348348 520774 348366
rect 491094 348268 520674 348348
rect 520754 348268 520774 348348
rect 491094 348230 520774 348268
rect 490953 348225 491099 348230
rect 490817 348096 490963 348101
rect 490817 347960 490822 348096
rect 490958 348062 520588 348096
rect 490958 347982 520454 348062
rect 520534 347982 520588 348062
rect 490958 347960 520588 347982
rect 490817 347955 490963 347960
rect 490817 347842 490963 347847
rect 490817 347706 490822 347842
rect 490958 347814 520410 347842
rect 490958 347734 520294 347814
rect 520374 347734 520410 347814
rect 490958 347706 520410 347734
rect 490817 347701 490963 347706
rect 490885 347572 491031 347577
rect 490885 347436 490890 347572
rect 491026 347548 520230 347572
rect 491026 347468 520134 347548
rect 520214 347468 520230 347548
rect 491026 347436 520230 347468
rect 490885 347431 491031 347436
rect 490935 347302 491081 347307
rect 490935 347166 490940 347302
rect 491076 347284 520094 347302
rect 491076 347204 519974 347284
rect 520054 347204 520094 347284
rect 491076 347166 520094 347204
rect 490935 347161 491081 347166
rect 452177 317803 453990 318107
rect 454294 317803 456177 318107
rect 452177 299098 456177 317803
rect 452177 292718 452458 299098
rect 455712 292718 456177 299098
rect 452177 278907 456177 292718
rect 452177 278603 453710 278907
rect 454014 278603 456177 278907
rect 452177 245525 456177 278603
rect 477612 283628 477920 283634
rect 477612 256611 477920 283320
rect 563796 261374 563802 261450
rect 563878 261374 563884 261450
rect 563802 260867 563878 261374
rect 563797 260862 563883 260867
rect 563797 260786 563802 260862
rect 563878 260786 563883 260862
rect 563797 260781 563883 260786
rect 563738 256972 563814 256978
rect 524989 256611 525307 256616
rect 477612 256303 524994 256611
rect 525302 256303 525307 256611
rect 563738 256519 563814 256896
rect 563733 256514 563819 256519
rect 563733 256438 563738 256514
rect 563814 256438 563819 256514
rect 563733 256433 563819 256438
rect 524989 256298 525307 256303
rect 563752 255436 563828 255442
rect 563752 254993 563828 255360
rect 563747 254988 563833 254993
rect 563747 254912 563752 254988
rect 563828 254912 563833 254988
rect 563747 254907 563833 254912
rect 524551 253331 524761 253336
rect 475878 253131 524556 253331
rect 524756 253131 524761 253331
rect 452177 245207 453947 245525
rect 454265 245207 456177 245525
rect 452177 205062 456177 245207
rect 452177 203816 453325 205062
rect 454571 203816 456177 205062
rect 452177 191899 456177 203816
rect 452177 187251 452333 191899
rect 455990 187251 456177 191899
rect 452177 177590 456177 187251
rect 452176 177478 456177 177590
rect 452176 176624 452276 177478
rect 456058 176624 456177 177478
rect 452176 176524 456177 176624
rect 444177 116216 445481 117462
rect 446727 116216 448177 117462
rect 444177 92247 448177 116216
rect 444177 91356 444290 92247
rect 448055 91356 448177 92247
rect 444177 74825 448177 91356
rect 444177 74534 446267 74825
rect 446558 74534 448177 74825
rect 436838 67677 437290 68598
rect 435826 67289 440158 67677
rect 159752 66158 162288 66334
rect 159752 63802 159964 66158
rect 162104 63802 162288 66158
rect 159752 63598 162288 63802
rect 435826 63691 436136 67289
rect 439734 63691 440158 67289
rect 435826 63345 440158 63691
rect 136832 58139 137772 59527
rect 139160 58139 140832 59527
rect 136832 43223 140832 58139
rect 444177 56044 448177 74534
rect 452177 115062 456177 176524
rect 452177 113816 453593 115062
rect 454839 113816 456177 115062
rect 452177 89388 456177 113816
rect 452177 88492 452241 89388
rect 456105 88492 456177 89388
rect 452177 73948 456177 88492
rect 452177 73571 453466 73948
rect 453843 73571 456177 73948
rect 452177 56044 456177 73571
rect 459575 246194 460533 246576
rect 475878 246194 476078 253131
rect 524551 253126 524761 253131
rect 524674 252974 525223 252979
rect 477763 252435 477769 252974
rect 478308 252435 524679 252974
rect 525218 252435 525223 252974
rect 524674 252430 525223 252435
rect 476829 247796 477147 247801
rect 459575 245994 476078 246194
rect 476828 247795 477148 247796
rect 476828 247477 476829 247795
rect 477147 247477 477148 247795
rect 136832 42905 138597 43223
rect 138915 42905 140832 43223
rect 136832 40865 140832 42905
rect 136832 31547 137083 40865
rect 140503 31547 140832 40865
rect 136832 30890 140832 31547
rect 3528 18157 4384 18189
rect 3528 17976 3562 18157
rect 1456 17822 3562 17976
rect 0 17710 1310 17822
rect 1430 17710 3562 17822
rect 1456 17563 3562 17710
rect 3528 17264 3562 17563
rect 4344 17264 4384 18157
rect 3528 17233 4384 17264
rect 124735 17233 124736 18189
rect 125692 17233 125693 18189
rect 124735 17232 125693 17233
rect 459575 18189 460533 245994
rect 476828 245526 477148 247477
rect 462580 245206 462586 245526
rect 462906 245206 477148 245526
rect 562634 244544 563019 244549
rect 462661 244169 462667 244544
rect 463042 244169 562639 244544
rect 563014 244169 563019 244544
rect 562634 244164 563019 244169
rect 564181 242632 564418 383151
rect 579257 382592 579494 471093
rect 580504 471076 580616 471082
rect 580504 455358 580616 470964
rect 583752 457058 583864 457064
rect 583752 456540 583864 456946
rect 583752 456428 584000 456540
rect 584112 456428 584800 456540
rect 580504 455246 584800 455358
rect 584320 454064 584800 454176
rect 584320 452882 584800 452994
rect 583194 451909 584160 451910
rect 583189 451647 583195 451909
rect 583457 451812 584160 451909
rect 583457 451700 585600 451812
rect 583457 451647 584160 451700
rect 583194 451646 584160 451647
rect 584320 450518 584800 450630
rect 583224 412118 583344 412126
rect 583224 412006 583228 412118
rect 583340 412006 583888 412118
rect 584000 412006 584800 412118
rect 583224 412000 583344 412006
rect 581531 410938 584447 410939
rect 581526 410854 581532 410938
rect 581616 410936 584447 410938
rect 581616 410854 584800 410936
rect 581531 410853 584800 410854
rect 584320 410824 584800 410853
rect 584320 409642 584800 409754
rect 584320 408460 584800 408572
rect 582282 407523 584160 407524
rect 582277 407261 582283 407523
rect 582545 407390 584160 407523
rect 582545 407278 585600 407390
rect 582545 407261 584160 407278
rect 582282 407260 584160 407261
rect 584320 406096 584800 406208
rect 531656 242396 564418 242632
rect 564859 382355 579494 382592
rect 531656 242395 563752 242396
rect 531656 185349 531893 242395
rect 564859 242148 565096 382355
rect 584320 365584 584800 365696
rect 584320 364480 584800 364514
rect 584288 364404 584800 364480
rect 584320 364402 584800 364404
rect 584320 363220 584800 363332
rect 584320 362038 584800 362150
rect 584320 360856 585600 360968
rect 584288 359674 584800 359786
rect 577993 356751 580972 356756
rect 577993 353782 577998 356751
rect 580967 353782 580972 356751
rect 577993 353777 580972 353782
rect 577998 349051 580967 353777
rect 577998 346076 580967 346082
rect 571755 319220 571976 323352
rect 570433 318999 571976 319220
rect 582226 320362 583886 320474
rect 583998 320362 585600 320474
rect 570433 311384 570654 318999
rect 571143 317802 571149 318108
rect 571455 317968 571855 318108
rect 582226 317968 582338 320362
rect 584178 319292 584444 319299
rect 584178 319268 585600 319292
rect 582954 319267 585600 319268
rect 582949 319193 582955 319267
rect 583029 319193 585600 319267
rect 582954 319192 585600 319193
rect 584178 319180 585600 319192
rect 584178 319179 584444 319180
rect 584320 317998 584800 318110
rect 571455 317856 582338 317968
rect 571455 317802 571855 317856
rect 571162 316872 571168 317192
rect 571488 316872 571912 317192
rect 584320 316816 584800 316928
rect 582511 315786 582773 315791
rect 582510 315785 584356 315786
rect 582510 315523 582511 315785
rect 582773 315747 584356 315785
rect 582773 315746 584383 315747
rect 582773 315634 584800 315746
rect 582773 315523 584356 315634
rect 582510 315522 584356 315523
rect 582511 315517 582773 315522
rect 584178 314452 585600 314564
rect 571048 311892 571054 312288
rect 571450 311892 572996 312288
rect 532234 241911 565096 242148
rect 565679 311163 570654 311384
rect 532234 185409 532471 241911
rect 565679 241632 565900 311163
rect 571062 310864 571068 311260
rect 571464 310864 571886 311260
rect 566898 310452 571738 310716
rect 582006 310452 582510 310716
rect 582774 310452 582780 310716
rect 532834 241411 565900 241632
rect 532834 185541 533055 241411
rect 566915 241116 567136 310452
rect 533414 240895 567136 241116
rect 531651 185114 531657 185349
rect 531892 185114 531898 185349
rect 532229 185174 532235 185409
rect 532470 185174 532476 185409
rect 532829 185322 532835 185541
rect 533054 185322 533060 185541
rect 532834 185321 533055 185322
rect 532234 185173 532471 185174
rect 531656 185113 531893 185114
rect 533414 179627 533635 240895
rect 570934 240343 571105 284149
rect 571461 278602 571467 278908
rect 571773 278820 571779 278908
rect 571773 278708 583920 278820
rect 571773 278602 571779 278708
rect 582686 276127 583490 276128
rect 582681 276053 582687 276127
rect 582761 276053 583490 276127
rect 582686 276052 583490 276053
rect 583566 276052 583572 276128
rect 583808 276052 583920 278708
rect 583808 275940 583996 276052
rect 584108 275940 585600 276052
rect 584112 274870 584437 274880
rect 584112 274858 585600 274870
rect 583252 274857 585600 274858
rect 583247 274783 583253 274857
rect 583327 274783 585600 274857
rect 583252 274782 585600 274783
rect 584112 274760 585600 274782
rect 584320 274758 585600 274760
rect 584320 273576 584800 273688
rect 571320 272692 571326 273088
rect 571722 272692 572996 273088
rect 584320 272394 584800 272506
rect 571276 271664 571282 272060
rect 571678 271664 571886 272060
rect 571258 271252 571738 271516
rect 582298 271368 583150 271516
rect 582298 271324 584436 271368
rect 582298 271252 584800 271324
rect 558218 240172 571105 240343
rect 533635 179406 534965 179584
rect 533414 179363 534965 179406
rect 558218 170466 558389 240172
rect 571261 239759 571387 271252
rect 582886 271212 584800 271252
rect 582886 271104 584436 271212
rect 584304 270030 585600 270142
rect 558751 239633 571387 239759
rect 574794 240690 584800 240830
rect 558213 170461 558394 170466
rect 558213 170290 558218 170461
rect 558389 170290 558394 170461
rect 558213 170285 558394 170290
rect 532226 161712 532234 161949
rect 532471 161712 534981 161949
rect 548989 151435 549292 151440
rect 510858 151142 510864 151435
rect 511157 151142 548994 151435
rect 549287 151142 549292 151435
rect 548989 151137 549292 151142
rect 549434 150748 549823 150753
rect 511035 150369 511041 150748
rect 511420 150369 549439 150748
rect 549818 150369 549823 150748
rect 549434 150364 549823 150369
rect 550001 149971 550675 155290
rect 510803 149297 510809 149971
rect 511483 149297 550675 149971
rect 511004 148158 511010 148778
rect 511630 148777 551648 148778
rect 511630 148159 551029 148777
rect 551647 148159 551653 148777
rect 511630 148158 551648 148159
rect 532828 81185 532834 81406
rect 533055 81185 536321 81406
rect 558751 73653 558877 239633
rect 574794 236252 574934 240690
rect 580058 236252 584800 240690
rect 574794 236030 584800 236252
rect 574794 230660 585600 230830
rect 574794 226222 574962 230660
rect 580086 226222 585600 230660
rect 574794 226030 585600 226222
rect 574794 196850 584800 197030
rect 574794 192412 574896 196850
rect 580020 192412 584800 196850
rect 574794 192230 584800 192412
rect 574794 186806 585600 187030
rect 574794 182368 574908 186806
rect 580032 182368 585600 186806
rect 574794 182230 585600 182368
rect 574794 152256 584800 152430
rect 574794 147818 575156 152256
rect 580280 147818 584800 152256
rect 574794 147630 584800 147818
rect 574794 142194 585600 142430
rect 574794 137756 575102 142194
rect 580226 137756 585600 142194
rect 574794 137630 585600 137756
rect 584320 96003 585600 96030
rect 584198 95929 585600 96003
rect 584320 95918 585600 95929
rect 584320 94818 585600 94848
rect 584198 94758 585600 94818
rect 584320 94736 585600 94758
rect 560528 93712 560747 93718
rect 560442 93554 560528 93666
rect 560747 93554 582624 93666
rect 584318 93554 584800 93666
rect 560528 93487 560747 93493
rect 582512 92484 582624 93554
rect 582512 92372 584076 92484
rect 584180 92372 584800 92484
rect 558746 73648 558882 73653
rect 558746 73522 558751 73648
rect 558877 73522 558882 73648
rect 558746 73517 558882 73522
rect 531650 63534 531656 63771
rect 531893 63534 536337 63771
rect 550541 55249 550844 55254
rect 527280 54956 527286 55249
rect 527579 54956 550546 55249
rect 550839 54956 550844 55249
rect 550541 54951 550844 54956
rect 527333 54732 527712 54738
rect 550986 54732 551375 54737
rect 527712 54353 550991 54732
rect 551370 54353 551375 54732
rect 527333 54347 527712 54353
rect 550986 54348 551375 54353
rect 551553 54009 552227 57112
rect 527689 53335 527695 54009
rect 528369 53335 552227 54009
rect 527846 52256 527852 52876
rect 528472 52875 553200 52876
rect 528472 52257 552581 52875
rect 553199 52257 553205 52875
rect 528472 52256 553200 52257
rect 584320 51344 585600 51372
rect 584196 51277 585600 51344
rect 584320 51260 585600 51277
rect 584320 50160 585600 50190
rect 583260 50091 585600 50160
rect 584320 50078 585600 50091
rect 532266 48896 532272 49008
rect 532384 48896 582642 49008
rect 584318 48896 584800 49008
rect 582530 47826 582642 48896
rect 582530 47714 583772 47826
rect 583894 47714 584800 47826
rect 584320 24878 585600 24914
rect 584304 24817 585600 24878
rect 584320 24802 585600 24817
rect 584320 23705 585600 23732
rect 583712 23644 585600 23705
rect 584320 23620 585600 23644
rect 532872 22438 532878 22550
rect 532990 22438 582906 22550
rect 584316 22438 584800 22550
rect 582794 21368 582906 22438
rect 582794 21256 583772 21368
rect 583898 21256 584800 21368
rect 584320 20142 585600 20186
rect 584216 20081 585600 20142
rect 584320 20074 585600 20081
rect 584320 18981 585600 19004
rect 583712 18920 585600 18981
rect 584320 18892 585600 18920
rect 459575 17233 459576 18189
rect 460532 17233 460533 18189
rect 531692 17710 531698 17822
rect 531810 17710 582690 17822
rect 584318 17710 584800 17822
rect 459575 17232 460533 17233
rect 124736 17227 125692 17232
rect 459576 17227 460532 17232
rect 582578 16640 582690 17710
rect 800 16528 1280 16640
rect 582578 16528 583488 16640
rect 583600 16528 584800 16640
rect 800 15346 1280 15458
rect 584320 15416 585600 15458
rect 584310 15355 585600 15416
rect 584320 15346 585600 15355
rect 448117 14678 448244 14683
rect 448117 14656 448122 14678
rect 448088 14576 448122 14656
rect 448117 14561 448122 14576
rect 448239 14656 448244 14678
rect 518029 14656 518119 14657
rect 448239 14652 518494 14656
rect 448239 14576 518034 14652
rect 448239 14561 448244 14576
rect 518029 14572 518034 14576
rect 518114 14576 518494 14652
rect 518114 14572 518119 14576
rect 518029 14567 518119 14572
rect 448117 14556 448244 14561
rect 450394 14491 518494 14496
rect 450394 14421 450515 14491
rect 450585 14488 518494 14491
rect 450585 14421 518194 14488
rect 450394 14416 518194 14421
rect 518189 14408 518194 14416
rect 518274 14416 518494 14488
rect 518274 14408 518279 14416
rect 518189 14403 518279 14408
rect 518349 14336 518439 14341
rect 451542 14331 518354 14336
rect 800 14164 1280 14276
rect 451542 14261 451699 14331
rect 451769 14261 518354 14331
rect 451542 14256 518354 14261
rect 518434 14256 518494 14336
rect 518349 14251 518439 14256
rect 584320 14241 585600 14276
rect 454044 14191 454144 14196
rect 454044 14176 454049 14191
rect 453978 14101 454049 14176
rect 454139 14176 454144 14191
rect 584294 14180 585600 14241
rect 518569 14176 518659 14179
rect 454139 14174 519190 14176
rect 454139 14101 518574 14174
rect 453978 14096 518574 14101
rect 518569 14094 518574 14096
rect 518654 14096 519190 14174
rect 584320 14164 585600 14180
rect 518654 14094 518659 14096
rect 518569 14089 518659 14094
rect 455228 14025 455328 14030
rect 455228 14016 455233 14025
rect 455148 13936 455233 14016
rect 455228 13935 455233 13936
rect 455323 14016 455328 14025
rect 518729 14022 518819 14027
rect 518729 14016 518734 14022
rect 455323 13942 518734 14016
rect 518814 14016 518819 14022
rect 518814 13942 519190 14016
rect 455323 13936 519190 13942
rect 455323 13935 455328 13936
rect 455228 13930 455328 13935
rect 457576 13857 457676 13862
rect 457576 13856 457581 13857
rect 457518 13776 457581 13856
rect 457576 13767 457581 13776
rect 457671 13856 457676 13857
rect 518889 13858 518979 13863
rect 518889 13856 518894 13858
rect 457671 13778 518894 13856
rect 518974 13856 518979 13858
rect 518974 13778 519190 13856
rect 457671 13776 519190 13778
rect 457671 13767 457676 13776
rect 518889 13773 518979 13776
rect 457576 13762 457676 13767
rect 458760 13699 458860 13704
rect 458760 13696 458765 13699
rect 458698 13616 458765 13696
rect 458760 13609 458765 13616
rect 458855 13696 458860 13699
rect 519049 13696 519139 13701
rect 458855 13616 519054 13696
rect 519134 13616 519190 13696
rect 458855 13609 458860 13616
rect 519049 13611 519139 13616
rect 458760 13604 458860 13609
rect 461127 13539 461227 13544
rect 461127 13536 461132 13539
rect 461100 13456 461132 13536
rect 76109 13450 76189 13452
rect 75554 13447 253278 13450
rect 75554 13377 76114 13447
rect 76184 13445 253278 13447
rect 76184 13377 253096 13445
rect 75554 13374 253096 13377
rect 253167 13374 253278 13445
rect 461127 13449 461132 13456
rect 461222 13536 461227 13539
rect 461222 13528 519898 13536
rect 461222 13456 519274 13528
rect 461222 13449 461227 13456
rect 461127 13444 461227 13449
rect 519269 13448 519274 13456
rect 519354 13456 519898 13528
rect 519354 13448 519359 13456
rect 519269 13443 519359 13448
rect 462311 13381 462411 13386
rect 462311 13376 462316 13381
rect 75554 13369 253278 13374
rect 462238 13296 462316 13376
rect 462311 13291 462316 13296
rect 462406 13376 462411 13381
rect 519429 13376 519519 13379
rect 462406 13374 519898 13376
rect 462406 13296 519434 13374
rect 462406 13291 462411 13296
rect 75554 13285 252090 13290
rect 462311 13286 462411 13291
rect 519429 13294 519434 13296
rect 519514 13296 519898 13374
rect 519514 13294 519519 13296
rect 519429 13289 519519 13294
rect 75554 13283 251904 13285
rect 75554 13213 75954 13283
rect 76024 13214 251904 13283
rect 251975 13214 252090 13285
rect 464671 13226 464765 13231
rect 464671 13216 464676 13226
rect 76024 13213 252090 13214
rect 75554 13209 252090 13213
rect 75949 13208 76029 13209
rect 464606 13142 464676 13216
rect 464760 13216 464765 13226
rect 519589 13216 519679 13221
rect 464760 13142 519594 13216
rect 464606 13136 519594 13142
rect 519674 13136 519898 13216
rect 519589 13131 519679 13136
rect 75554 13125 249712 13130
rect 75554 13121 249554 13125
rect 0 12982 1280 13094
rect 75554 13051 75794 13121
rect 75864 13054 249554 13121
rect 249625 13054 249712 13125
rect 465855 13060 465949 13065
rect 465855 13056 465860 13060
rect 75864 13051 249712 13054
rect 75554 13049 249712 13051
rect 75789 13046 75869 13049
rect 465770 12976 465860 13056
rect 465944 13056 465949 13060
rect 519749 13056 519839 13061
rect 465944 12976 519754 13056
rect 519834 12976 519898 13056
rect 584320 12982 584800 13094
rect 465855 12971 465949 12976
rect 519749 12971 519839 12976
rect 75554 12965 248508 12970
rect 75554 12963 248370 12965
rect 75554 12893 75634 12963
rect 75704 12894 248370 12963
rect 248441 12894 248508 12965
rect 468222 12896 468316 12899
rect 519969 12898 520059 12903
rect 519969 12896 519974 12898
rect 75704 12893 248508 12894
rect 75554 12889 248508 12893
rect 468154 12894 519974 12896
rect 75629 12888 75709 12889
rect 468154 12816 468227 12894
rect 246006 12811 246106 12816
rect 246006 12810 246011 12811
rect 74850 12803 246011 12810
rect 74850 12733 75414 12803
rect 75484 12733 246011 12803
rect 74850 12729 246011 12733
rect 75409 12728 75489 12729
rect 246006 12721 246011 12729
rect 246101 12810 246106 12811
rect 468222 12810 468227 12816
rect 468311 12818 519974 12894
rect 520054 12896 520059 12898
rect 520054 12818 520608 12896
rect 468311 12816 520608 12818
rect 468311 12810 468316 12816
rect 519969 12813 520059 12816
rect 246101 12729 246134 12810
rect 468222 12805 468316 12810
rect 469406 12738 469500 12743
rect 469406 12736 469411 12738
rect 246101 12721 246106 12729
rect 246006 12716 246106 12721
rect 469326 12656 469411 12736
rect 244822 12651 244922 12656
rect 244822 12650 244827 12651
rect 74850 12643 244827 12650
rect 74850 12573 75254 12643
rect 75324 12573 244827 12643
rect 74850 12569 244827 12573
rect 75249 12568 75329 12569
rect 244822 12561 244827 12569
rect 244917 12650 244922 12651
rect 469406 12654 469411 12656
rect 469495 12736 469500 12738
rect 520129 12738 520219 12743
rect 520129 12736 520134 12738
rect 469495 12658 520134 12736
rect 520214 12736 520219 12738
rect 520214 12658 520608 12736
rect 469495 12656 520608 12658
rect 469495 12654 469500 12656
rect 244917 12569 244946 12650
rect 469406 12649 469500 12654
rect 520129 12653 520219 12656
rect 471763 12576 471857 12579
rect 520289 12578 520379 12583
rect 520289 12576 520294 12578
rect 471704 12574 520294 12576
rect 244917 12561 244922 12569
rect 244822 12556 244922 12561
rect 242470 12497 242570 12502
rect 242470 12490 242475 12497
rect 74850 12481 242475 12490
rect 74850 12411 75094 12481
rect 75164 12411 242475 12481
rect 74850 12409 242475 12411
rect 75089 12406 75169 12409
rect 242470 12407 242475 12409
rect 242565 12490 242570 12497
rect 471704 12496 471768 12574
rect 471763 12490 471768 12496
rect 471852 12498 520294 12574
rect 520374 12576 520379 12578
rect 520374 12498 520608 12576
rect 471852 12496 520608 12498
rect 471852 12490 471857 12496
rect 520289 12493 520379 12496
rect 242565 12409 242606 12490
rect 471763 12485 471857 12490
rect 472947 12416 473041 12419
rect 520449 12418 520539 12423
rect 520449 12416 520454 12418
rect 472892 12414 520454 12416
rect 242565 12407 242570 12409
rect 242470 12402 242570 12407
rect 241286 12335 241386 12340
rect 472892 12336 472952 12414
rect 241286 12330 241291 12335
rect 74850 12325 241291 12330
rect 74850 12255 74934 12325
rect 75004 12255 241291 12325
rect 74850 12249 241291 12255
rect 241286 12245 241291 12249
rect 241381 12330 241386 12335
rect 472947 12330 472952 12336
rect 473036 12338 520454 12414
rect 520534 12416 520539 12418
rect 520534 12338 520608 12416
rect 473036 12336 520608 12338
rect 473036 12330 473041 12336
rect 520449 12333 520539 12336
rect 241381 12249 241408 12330
rect 472947 12325 473041 12330
rect 475314 12264 475408 12269
rect 475314 12256 475319 12264
rect 241381 12245 241386 12249
rect 241286 12240 241386 12245
rect 475236 12180 475319 12256
rect 475403 12256 475408 12264
rect 520669 12256 520759 12261
rect 475403 12180 520674 12256
rect 238922 12173 239022 12178
rect 475236 12176 520674 12180
rect 520754 12176 521278 12256
rect 475314 12175 475408 12176
rect 238922 12170 238927 12173
rect 74146 12161 238927 12170
rect 74146 12091 74714 12161
rect 74784 12091 238927 12161
rect 74146 12089 238927 12091
rect 74709 12086 74789 12089
rect 238922 12083 238927 12089
rect 239017 12170 239022 12173
rect 520669 12171 520759 12176
rect 239017 12089 239054 12170
rect 476498 12100 476592 12105
rect 476498 12096 476503 12100
rect 239017 12083 239022 12089
rect 238922 12078 239022 12083
rect 476406 12016 476503 12096
rect 476587 12096 476592 12100
rect 520829 12098 520919 12103
rect 520829 12096 520834 12098
rect 476587 12018 520834 12096
rect 520914 12096 520919 12098
rect 520914 12018 521278 12096
rect 476587 12016 521278 12018
rect 237738 12011 237838 12016
rect 476498 12011 476592 12016
rect 520829 12013 520919 12016
rect 237738 12010 237743 12011
rect 74146 12003 237743 12010
rect 74146 11933 74554 12003
rect 74624 11933 237743 12003
rect 74146 11929 237743 11933
rect 74549 11928 74629 11929
rect 237738 11921 237743 11929
rect 237833 12010 237838 12011
rect 237833 11929 237872 12010
rect 478864 11940 478958 11945
rect 478864 11936 478869 11940
rect 237833 11921 237838 11929
rect 237738 11916 237838 11921
rect 0 11800 1280 11912
rect 235357 11854 235467 11859
rect 478800 11856 478869 11936
rect 478953 11936 478958 11940
rect 520989 11936 521079 11941
rect 478953 11856 520994 11936
rect 521074 11856 521278 11936
rect 235357 11850 235362 11854
rect 74146 11845 235362 11850
rect 74146 11775 74394 11845
rect 74464 11775 235362 11845
rect 74146 11769 235362 11775
rect 235357 11754 235362 11769
rect 235462 11850 235467 11854
rect 478864 11851 478958 11856
rect 520989 11851 521079 11856
rect 235462 11769 235480 11850
rect 584320 11800 584800 11912
rect 480048 11782 480142 11787
rect 480048 11776 480053 11782
rect 235462 11754 235467 11769
rect 235357 11749 235467 11754
rect 234173 11696 234283 11701
rect 479998 11698 480053 11776
rect 480137 11776 480142 11782
rect 521149 11776 521239 11781
rect 480137 11698 521154 11776
rect 479998 11696 521154 11698
rect 521234 11696 521278 11776
rect 234173 11690 234178 11696
rect 74146 11681 234178 11690
rect 74146 11611 74234 11681
rect 74304 11611 234178 11681
rect 74146 11609 234178 11611
rect 74229 11606 74309 11609
rect 234173 11596 234178 11609
rect 234278 11690 234283 11696
rect 480048 11693 480142 11696
rect 521149 11691 521239 11696
rect 234278 11609 234294 11690
rect 482410 11621 482495 11626
rect 482410 11616 482415 11621
rect 234278 11596 234283 11609
rect 234173 11591 234283 11596
rect 231809 11542 231919 11547
rect 231809 11530 231814 11542
rect 73444 11523 231814 11530
rect 73444 11453 74014 11523
rect 74084 11453 231814 11523
rect 73444 11449 231814 11453
rect 74009 11448 74089 11449
rect 231809 11442 231814 11449
rect 231914 11530 231919 11542
rect 482316 11546 482415 11616
rect 482490 11616 482495 11621
rect 521369 11616 521459 11619
rect 482490 11614 521988 11616
rect 482490 11546 521374 11614
rect 482316 11536 521374 11546
rect 521369 11534 521374 11536
rect 521454 11536 521988 11614
rect 521454 11534 521459 11536
rect 231914 11449 231976 11530
rect 521369 11529 521459 11534
rect 483594 11456 483679 11460
rect 521529 11458 521619 11463
rect 521529 11456 521534 11458
rect 483530 11455 521534 11456
rect 231914 11442 231919 11449
rect 231809 11437 231919 11442
rect 230625 11384 230735 11389
rect 230625 11370 230630 11384
rect 73444 11363 230630 11370
rect 73444 11293 73854 11363
rect 73924 11293 230630 11363
rect 73444 11289 230630 11293
rect 73849 11288 73929 11289
rect 230625 11284 230630 11289
rect 230730 11370 230735 11384
rect 483530 11380 483599 11455
rect 483674 11380 521534 11455
rect 483530 11378 521534 11380
rect 521614 11456 521619 11458
rect 521614 11378 521988 11456
rect 483530 11376 521988 11378
rect 483594 11375 483679 11376
rect 521529 11373 521619 11376
rect 230730 11289 230758 11370
rect 485951 11299 486036 11304
rect 485951 11296 485956 11299
rect 230730 11284 230735 11289
rect 230625 11279 230735 11284
rect 228283 11224 228393 11229
rect 228283 11210 228288 11224
rect 73444 11201 228288 11210
rect 73444 11131 73694 11201
rect 73764 11131 228288 11201
rect 73444 11129 228288 11131
rect 73689 11126 73769 11129
rect 228283 11124 228288 11129
rect 228388 11210 228393 11224
rect 485890 11224 485956 11296
rect 486031 11296 486036 11299
rect 486031 11288 521988 11296
rect 486031 11224 521694 11288
rect 485890 11216 521694 11224
rect 228388 11129 228440 11210
rect 521689 11208 521694 11216
rect 521774 11216 521988 11288
rect 521774 11208 521779 11216
rect 521689 11203 521779 11208
rect 487135 11139 487220 11144
rect 487135 11136 487140 11139
rect 228388 11124 228393 11129
rect 228283 11119 228393 11124
rect 227099 11060 227209 11065
rect 73529 11050 73609 11052
rect 227099 11050 227104 11060
rect 73444 11047 227104 11050
rect 73444 10977 73534 11047
rect 73604 10977 227104 11047
rect 73444 10969 227104 10977
rect 227099 10960 227104 10969
rect 227204 11050 227209 11060
rect 487052 11064 487140 11136
rect 487215 11136 487220 11139
rect 521849 11136 521939 11141
rect 487215 11064 521854 11136
rect 487052 11056 521854 11064
rect 521934 11056 521988 11136
rect 521849 11051 521939 11056
rect 227204 10969 227248 11050
rect 489473 10976 489558 10978
rect 522069 10976 522159 10979
rect 489388 10974 522696 10976
rect 489388 10973 522074 10974
rect 227204 10960 227209 10969
rect 227099 10955 227209 10960
rect 224735 10900 224845 10905
rect 224735 10890 224740 10900
rect 72730 10883 224740 10890
rect 72730 10813 73314 10883
rect 73384 10813 224740 10883
rect 72730 10809 224740 10813
rect 73309 10808 73389 10809
rect 224735 10800 224740 10809
rect 224840 10890 224845 10900
rect 489388 10898 489478 10973
rect 489553 10898 522074 10973
rect 489388 10896 522074 10898
rect 489473 10893 489558 10896
rect 522069 10894 522074 10896
rect 522154 10896 522696 10974
rect 522154 10894 522159 10896
rect 224840 10809 224892 10890
rect 522069 10889 522159 10894
rect 490657 10817 490742 10822
rect 490657 10816 490662 10817
rect 224840 10800 224845 10809
rect 224735 10795 224845 10800
rect 223551 10742 223661 10747
rect 223551 10730 223556 10742
rect 800 10618 1280 10730
rect 72730 10723 223556 10730
rect 72730 10653 73154 10723
rect 73224 10653 223556 10723
rect 72730 10649 223556 10653
rect 73149 10648 73229 10649
rect 223551 10642 223556 10649
rect 223656 10730 223661 10742
rect 490592 10742 490662 10816
rect 490737 10816 490742 10817
rect 490737 10810 522696 10816
rect 490737 10742 522234 10810
rect 490592 10736 522234 10742
rect 522229 10730 522234 10736
rect 522314 10736 522696 10810
rect 522314 10730 522319 10736
rect 223656 10649 223692 10730
rect 522229 10725 522319 10730
rect 584320 10716 585600 10730
rect 493043 10656 493128 10660
rect 522389 10656 522479 10657
rect 492970 10655 522696 10656
rect 223656 10642 223661 10649
rect 223551 10637 223661 10642
rect 221197 10584 221307 10589
rect 221197 10570 221202 10584
rect 72730 10565 221202 10570
rect 72730 10495 72994 10565
rect 73064 10495 221202 10565
rect 72730 10489 221202 10495
rect 221197 10484 221202 10489
rect 221302 10570 221307 10584
rect 492970 10580 493048 10655
rect 493123 10652 522696 10655
rect 493123 10580 522394 10652
rect 492970 10576 522394 10580
rect 493043 10575 493128 10576
rect 221302 10489 221322 10570
rect 294481 10568 294551 10573
rect 522389 10572 522394 10576
rect 522474 10576 522696 10652
rect 584276 10635 585600 10716
rect 584320 10618 585600 10635
rect 522474 10572 522479 10576
rect 282622 10544 294486 10568
rect 221302 10484 221307 10489
rect 282622 10488 282707 10544
rect 221197 10479 221307 10484
rect 282702 10484 282707 10488
rect 282767 10508 294486 10544
rect 294546 10508 294648 10568
rect 522389 10567 522479 10572
rect 282767 10488 294648 10508
rect 494227 10499 494312 10504
rect 494227 10496 494232 10499
rect 282767 10484 282772 10488
rect 282702 10479 282772 10484
rect 220013 10422 220123 10427
rect 220013 10410 220018 10422
rect 72730 10405 220018 10410
rect 72730 10335 72834 10405
rect 72904 10335 220018 10405
rect 72730 10329 220018 10335
rect 220013 10322 220018 10329
rect 220118 10410 220123 10422
rect 494134 10424 494232 10496
rect 494307 10496 494312 10499
rect 522549 10496 522639 10499
rect 494307 10494 522696 10496
rect 494307 10424 522554 10494
rect 494134 10416 522554 10424
rect 220118 10329 220178 10410
rect 282422 10408 282492 10411
rect 290933 10410 291003 10415
rect 290933 10408 290938 10410
rect 282332 10406 290938 10408
rect 282332 10346 282427 10406
rect 282487 10350 290938 10406
rect 290998 10408 291003 10410
rect 522549 10414 522554 10416
rect 522634 10416 522696 10494
rect 522634 10414 522639 10416
rect 522549 10409 522639 10414
rect 290998 10350 291112 10408
rect 282487 10346 291112 10350
rect 220118 10322 220123 10329
rect 282332 10328 291112 10346
rect 522769 10336 522859 10337
rect 496494 10332 523368 10336
rect 220013 10317 220123 10322
rect 496494 10327 522774 10332
rect 287386 10252 287456 10257
rect 496494 10256 496589 10327
rect 72036 10245 217782 10250
rect 287386 10248 287391 10252
rect 72036 10243 217658 10245
rect 72036 10173 72614 10243
rect 72684 10174 217658 10243
rect 217729 10174 217782 10245
rect 72684 10173 217782 10174
rect 72036 10169 217782 10173
rect 282042 10228 287391 10248
rect 72609 10168 72689 10169
rect 282042 10168 282147 10228
rect 282207 10192 287391 10228
rect 287451 10248 287456 10252
rect 496584 10252 496589 10256
rect 496664 10256 522774 10327
rect 496664 10252 496669 10256
rect 287451 10192 287530 10248
rect 496584 10247 496669 10252
rect 522769 10252 522774 10256
rect 522854 10256 523368 10332
rect 522854 10252 522859 10256
rect 522769 10247 522859 10252
rect 282207 10168 287530 10192
rect 522929 10178 523019 10183
rect 522929 10176 522934 10178
rect 497674 10171 522934 10176
rect 282142 10163 282212 10168
rect 283838 10102 283908 10107
rect 72036 10085 216600 10090
rect 283838 10088 283843 10102
rect 72036 10015 72454 10085
rect 72524 10015 216476 10085
rect 72036 10014 216476 10015
rect 216547 10014 216600 10085
rect 72036 10009 216600 10014
rect 281786 10066 283843 10088
rect 281786 10008 281867 10066
rect 281862 10006 281867 10008
rect 281927 10042 283843 10066
rect 283903 10088 283908 10102
rect 497674 10096 497773 10171
rect 497848 10098 522934 10171
rect 523014 10176 523019 10178
rect 523014 10098 523368 10176
rect 497848 10096 523368 10098
rect 497768 10091 497853 10096
rect 522929 10093 523019 10096
rect 283903 10042 283974 10088
rect 281927 10008 283974 10042
rect 523089 10026 523179 10031
rect 500135 10016 500220 10020
rect 523089 10016 523094 10026
rect 500068 10015 523094 10016
rect 281927 10006 281932 10008
rect 281862 10001 281932 10006
rect 280291 9936 280361 9941
rect 500068 9940 500140 10015
rect 500215 9946 523094 10015
rect 523174 10016 523179 10026
rect 523174 9946 523368 10016
rect 500215 9940 523368 9946
rect 500068 9936 523368 9940
rect 72036 9925 214290 9930
rect 280291 9928 280296 9936
rect 72036 9855 72294 9925
rect 72364 9920 214290 9925
rect 72364 9855 214129 9920
rect 72036 9851 214129 9855
rect 214198 9851 214290 9920
rect 72036 9849 214290 9851
rect 280196 9876 280296 9928
rect 280356 9928 280361 9936
rect 500135 9935 500220 9936
rect 280356 9912 281702 9928
rect 280356 9876 281587 9912
rect 280196 9852 281587 9876
rect 281647 9852 281702 9912
rect 523249 9856 523339 9857
rect 214124 9846 214203 9849
rect 280196 9848 281702 9852
rect 501282 9852 523368 9856
rect 501282 9851 523254 9852
rect 281582 9847 281652 9848
rect 501282 9776 501324 9851
rect 501399 9776 523254 9851
rect 501319 9771 501404 9776
rect 523249 9772 523254 9776
rect 523334 9776 523368 9852
rect 523334 9772 523339 9776
rect 72036 9765 213078 9770
rect 72036 9695 72134 9765
rect 72204 9758 213078 9765
rect 72204 9695 212945 9758
rect 72036 9689 212945 9695
rect 213014 9689 213078 9758
rect 276658 9760 281448 9768
rect 523249 9767 523339 9772
rect 276658 9700 276749 9760
rect 276809 9750 281448 9760
rect 276809 9700 281307 9750
rect 276658 9690 281307 9700
rect 281367 9690 281448 9750
rect 212940 9684 213019 9689
rect 276658 9688 281448 9690
rect 503624 9690 524100 9696
rect 281302 9685 281372 9688
rect 503624 9684 523474 9690
rect 503624 9624 503689 9684
rect 503749 9624 523474 9684
rect 503624 9616 523474 9624
rect 71909 9610 71989 9612
rect 273196 9610 273266 9615
rect 71390 9607 210696 9610
rect 273196 9608 273201 9610
rect 800 9543 42536 9548
rect 800 9441 42429 9543
rect 42531 9441 42536 9543
rect 71390 9537 71914 9607
rect 71984 9596 210696 9607
rect 71984 9537 210577 9596
rect 71390 9529 210577 9537
rect 210572 9527 210577 9529
rect 210646 9529 210696 9596
rect 273152 9550 273201 9608
rect 273261 9608 273266 9610
rect 523469 9610 523474 9616
rect 523554 9616 524100 9690
rect 523554 9610 523559 9616
rect 273261 9588 281142 9608
rect 523469 9605 523559 9610
rect 273261 9550 281027 9588
rect 210646 9527 210651 9529
rect 273152 9528 281027 9550
rect 281087 9528 281142 9588
rect 523629 9538 523719 9543
rect 523629 9536 523634 9538
rect 210572 9522 210651 9527
rect 281022 9523 281092 9528
rect 504788 9524 523634 9536
rect 504788 9464 504873 9524
rect 504933 9464 523634 9524
rect 504788 9458 523634 9464
rect 523714 9536 523719 9538
rect 523714 9458 524100 9536
rect 584320 9530 585600 9548
rect 584300 9463 585600 9530
rect 504788 9456 524100 9458
rect 523629 9453 523719 9456
rect 800 9436 42536 9441
rect 71390 9445 209526 9450
rect 71390 9375 71754 9445
rect 71824 9438 209526 9445
rect 71824 9375 209393 9438
rect 71390 9369 209393 9375
rect 209462 9369 209526 9438
rect 297940 9442 304098 9448
rect 297940 9440 303962 9442
rect 297940 9380 298033 9440
rect 298093 9382 303962 9440
rect 304022 9382 304098 9442
rect 584320 9436 585600 9463
rect 298093 9380 304098 9382
rect 209388 9364 209467 9369
rect 297940 9368 304098 9380
rect 507198 9370 524100 9376
rect 507198 9368 523794 9370
rect 507198 9308 507249 9368
rect 507309 9308 523794 9368
rect 207014 9292 207093 9297
rect 507198 9296 523794 9308
rect 207014 9290 207019 9292
rect 71390 9285 207019 9290
rect 71390 9215 71594 9285
rect 71664 9223 207019 9285
rect 207088 9290 207093 9292
rect 523789 9290 523794 9296
rect 523874 9296 524100 9370
rect 523874 9290 523879 9296
rect 207088 9223 207138 9290
rect 71664 9215 207138 9223
rect 71390 9209 207138 9215
rect 301468 9282 304430 9288
rect 523789 9285 523879 9290
rect 301468 9222 301569 9282
rect 301629 9272 304430 9282
rect 301629 9222 304242 9272
rect 301468 9212 304242 9222
rect 304302 9212 304430 9272
rect 508428 9216 508498 9221
rect 523949 9216 524039 9221
rect 301468 9208 304430 9212
rect 304237 9207 304307 9208
rect 508354 9156 508433 9216
rect 508493 9156 523954 9216
rect 6258 9147 42850 9152
rect 6258 9045 42743 9147
rect 42845 9045 42850 9147
rect 205830 9134 205909 9139
rect 508354 9136 523954 9156
rect 524034 9136 524100 9216
rect 205830 9130 205835 9134
rect 71390 9121 205835 9130
rect 71390 9051 71434 9121
rect 71504 9065 205835 9121
rect 205904 9130 205909 9134
rect 205904 9065 206002 9130
rect 306117 9128 306187 9133
rect 523949 9131 524039 9136
rect 71504 9051 206002 9065
rect 71390 9049 206002 9051
rect 304412 9118 306122 9128
rect 304412 9058 304522 9118
rect 304582 9068 306122 9118
rect 306182 9068 306228 9128
rect 304582 9058 306228 9068
rect 71429 9046 71509 9049
rect 304412 9048 306228 9058
rect 524169 9056 524259 9059
rect 510714 9054 524808 9056
rect 510714 9046 524174 9054
rect 6258 9040 42850 9045
rect 0 8254 1280 8366
rect 0 7072 1280 7184
rect 800 5890 1280 6002
rect 6258 4820 6370 9040
rect 510714 8986 510800 9046
rect 510860 8986 524174 9046
rect 510714 8976 524174 8986
rect 524169 8974 524174 8976
rect 524254 8976 524808 9054
rect 524254 8974 524259 8976
rect 70686 8963 203632 8970
rect 524169 8969 524259 8974
rect 70686 8893 71214 8963
rect 71284 8960 203632 8963
rect 71284 8900 203478 8960
rect 203538 8900 203632 8960
rect 71284 8893 203632 8900
rect 70686 8889 203632 8893
rect 304734 8962 308874 8968
rect 304734 8956 308682 8962
rect 304734 8896 304802 8956
rect 304862 8902 308682 8956
rect 308742 8902 308874 8962
rect 304862 8896 308874 8902
rect 524329 8896 524419 8901
rect 71209 8888 71289 8889
rect 304734 8888 308874 8896
rect 511918 8886 524334 8896
rect 511918 8826 511984 8886
rect 512044 8826 524334 8886
rect 511918 8816 524334 8826
rect 524414 8816 524808 8896
rect 312205 8810 312275 8815
rect 524329 8811 524419 8816
rect 70686 8803 202446 8810
rect 312205 8808 312210 8810
rect 70686 8733 71054 8803
rect 71124 8802 202446 8803
rect 71124 8742 202294 8802
rect 202354 8742 202446 8802
rect 71124 8733 202446 8742
rect 70686 8729 202446 8733
rect 305040 8778 312210 8808
rect 71049 8728 71129 8729
rect 305040 8728 305082 8778
rect 305077 8718 305082 8728
rect 305142 8750 312210 8778
rect 312270 8808 312275 8810
rect 312270 8750 312328 8808
rect 305142 8728 312328 8750
rect 524489 8738 524579 8743
rect 524489 8736 524494 8738
rect 514262 8730 524494 8736
rect 305142 8718 305147 8728
rect 305077 8713 305147 8718
rect 199915 8661 200015 8666
rect 199915 8650 199920 8661
rect 70686 8643 199920 8650
rect 70686 8573 70894 8643
rect 70964 8573 199920 8643
rect 70686 8571 199920 8573
rect 200010 8650 200015 8661
rect 315765 8660 315835 8665
rect 200010 8571 200062 8650
rect 315765 8648 315770 8660
rect 70686 8569 200062 8571
rect 305328 8632 315770 8648
rect 305328 8572 305362 8632
rect 305422 8600 315770 8632
rect 315830 8648 315835 8660
rect 514262 8656 514324 8730
rect 514319 8654 514324 8656
rect 514400 8658 524494 8730
rect 524574 8736 524579 8738
rect 524574 8658 524808 8736
rect 514400 8656 524808 8658
rect 514400 8654 514405 8656
rect 514319 8649 514405 8654
rect 524489 8653 524579 8656
rect 315830 8600 315924 8648
rect 305422 8572 315924 8600
rect 70889 8568 70969 8569
rect 199915 8566 200015 8569
rect 305328 8568 315924 8572
rect 515442 8570 524808 8576
rect 305357 8567 305427 8568
rect 515442 8496 515508 8570
rect 198731 8491 198831 8496
rect 515503 8494 515508 8496
rect 515584 8496 524654 8570
rect 515584 8494 515589 8496
rect 198731 8490 198736 8491
rect 70686 8483 198736 8490
rect 70686 8413 70734 8483
rect 70804 8413 198736 8483
rect 70686 8409 198736 8413
rect 70729 8408 70809 8409
rect 198731 8401 198736 8409
rect 198826 8490 198831 8491
rect 198826 8409 198862 8490
rect 305637 8488 305707 8491
rect 515503 8489 515589 8494
rect 524649 8490 524654 8496
rect 524734 8496 524808 8570
rect 524734 8490 524739 8496
rect 319304 8488 319374 8489
rect 305592 8486 319478 8488
rect 305592 8426 305642 8486
rect 305702 8484 319478 8486
rect 524649 8485 524739 8490
rect 305702 8426 319309 8484
rect 305592 8424 319309 8426
rect 319369 8424 319478 8484
rect 198826 8401 198831 8409
rect 305592 8408 319478 8424
rect 517869 8416 517955 8419
rect 524869 8416 524959 8419
rect 517776 8414 525468 8416
rect 198731 8396 198831 8401
rect 196354 8339 196454 8344
rect 196354 8330 196359 8339
rect 21658 8323 196359 8330
rect 21658 8253 22214 8323
rect 22284 8253 196359 8323
rect 21658 8249 196359 8253
rect 196449 8330 196454 8339
rect 517776 8338 517874 8414
rect 517950 8338 524874 8414
rect 517776 8336 524874 8338
rect 517869 8333 517955 8336
rect 524869 8334 524874 8336
rect 524954 8336 525468 8414
rect 524954 8334 524959 8336
rect 196449 8249 196520 8330
rect 524869 8329 524959 8334
rect 525029 8260 525119 8265
rect 519053 8256 519139 8259
rect 525029 8256 525034 8260
rect 518974 8254 525034 8256
rect 22209 8248 22289 8249
rect 196354 8244 196454 8249
rect 518974 8178 519058 8254
rect 519134 8180 525034 8254
rect 525114 8256 525119 8260
rect 525114 8180 525468 8256
rect 584320 8254 584800 8366
rect 519134 8178 525468 8180
rect 195170 8173 195270 8178
rect 518974 8176 525468 8178
rect 519053 8173 519139 8176
rect 525029 8175 525119 8176
rect 22049 8170 22129 8172
rect 195170 8170 195175 8173
rect 21658 8167 195175 8170
rect 21658 8097 22054 8167
rect 22124 8097 195175 8167
rect 21658 8089 195175 8097
rect 195170 8083 195175 8089
rect 195265 8170 195270 8173
rect 195265 8089 195320 8170
rect 525189 8096 525279 8101
rect 521334 8090 525194 8096
rect 195265 8083 195270 8089
rect 195170 8078 195270 8083
rect 521334 8016 521425 8090
rect 521420 8014 521425 8016
rect 521501 8016 525194 8090
rect 525274 8016 525468 8096
rect 521501 8014 521506 8016
rect 21658 8005 192944 8010
rect 521420 8009 521506 8014
rect 525189 8011 525279 8016
rect 21658 7935 21894 8005
rect 21964 7991 192944 8005
rect 21964 7935 192827 7991
rect 21658 7929 192827 7935
rect 192822 7921 192827 7929
rect 192897 7929 192944 7991
rect 539349 7940 539439 7945
rect 539349 7936 539354 7940
rect 522522 7930 539354 7936
rect 192897 7921 192902 7929
rect 192822 7916 192902 7921
rect 522522 7856 522609 7930
rect 522604 7854 522609 7856
rect 522685 7860 539354 7930
rect 539434 7936 539439 7940
rect 539434 7860 539468 7936
rect 522685 7856 539468 7860
rect 522685 7854 522690 7856
rect 539349 7855 539439 7856
rect 191638 7850 191718 7854
rect 21658 7849 191770 7850
rect 522604 7849 522690 7854
rect 21658 7845 191643 7849
rect 21658 7775 21734 7845
rect 21804 7779 191643 7845
rect 191713 7779 191770 7849
rect 21804 7775 191770 7779
rect 539569 7778 539659 7783
rect 524971 7776 525057 7777
rect 539569 7776 539574 7778
rect 21658 7769 191770 7775
rect 524950 7772 539574 7776
rect 189282 7694 189373 7699
rect 524950 7696 524976 7772
rect 525052 7698 539574 7772
rect 539654 7776 539659 7778
rect 539654 7698 540176 7776
rect 525052 7696 540176 7698
rect 189282 7690 189287 7694
rect 20632 7683 189287 7690
rect 20632 7613 21214 7683
rect 21284 7613 189287 7683
rect 189368 7690 189373 7694
rect 524971 7691 525057 7696
rect 539569 7693 539659 7696
rect 189368 7613 189404 7690
rect 539729 7624 539819 7629
rect 526155 7616 526241 7621
rect 539729 7616 539734 7624
rect 20632 7609 189404 7613
rect 21209 7608 21289 7609
rect 189282 7608 189373 7609
rect 526138 7540 526160 7616
rect 526236 7544 539734 7616
rect 539814 7616 539819 7624
rect 539814 7544 540176 7616
rect 526236 7540 540176 7544
rect 526138 7536 540176 7540
rect 526155 7535 526241 7536
rect 20632 7521 188218 7530
rect 20632 7451 21054 7521
rect 21124 7520 188218 7521
rect 21124 7451 188103 7520
rect 20632 7449 188103 7451
rect 21049 7446 21129 7449
rect 188098 7439 188103 7449
rect 188184 7449 188218 7520
rect 539889 7466 539979 7471
rect 528503 7458 528589 7463
rect 528503 7456 528508 7458
rect 188184 7439 188189 7449
rect 188098 7434 188189 7439
rect 528478 7382 528508 7456
rect 528584 7456 528589 7458
rect 539889 7456 539894 7466
rect 528584 7386 539894 7456
rect 539974 7456 539979 7466
rect 539974 7386 540176 7456
rect 528584 7382 540176 7386
rect 185742 7372 185833 7377
rect 528478 7376 540176 7382
rect 185742 7370 185747 7372
rect 20632 7361 185747 7370
rect 20632 7291 20894 7361
rect 20964 7291 185747 7361
rect 185828 7370 185833 7372
rect 185828 7291 185882 7370
rect 529687 7302 529773 7307
rect 529687 7296 529692 7302
rect 20632 7289 185882 7291
rect 20889 7286 20969 7289
rect 185742 7286 185833 7289
rect 529586 7226 529692 7296
rect 529768 7296 529773 7302
rect 540049 7296 540139 7299
rect 529768 7294 540176 7296
rect 529768 7226 540054 7294
rect 184558 7218 184649 7223
rect 184558 7210 184563 7218
rect 20632 7203 184563 7210
rect 20632 7133 20734 7203
rect 20804 7137 184563 7203
rect 184644 7210 184649 7218
rect 529586 7216 540054 7226
rect 540049 7214 540054 7216
rect 540134 7216 540176 7294
rect 540134 7214 540139 7216
rect 184644 7137 184712 7210
rect 540049 7209 540139 7214
rect 20804 7133 184712 7137
rect 532044 7142 532130 7147
rect 532044 7136 532049 7142
rect 20632 7129 184712 7133
rect 20729 7128 20809 7129
rect 531972 7066 532049 7136
rect 532125 7136 532130 7142
rect 540269 7142 540359 7147
rect 540269 7136 540274 7142
rect 532125 7066 540274 7136
rect 531972 7062 540274 7066
rect 540354 7136 540359 7142
rect 540354 7062 540896 7136
rect 584320 7072 584800 7184
rect 531972 7056 540896 7062
rect 182178 7050 182269 7055
rect 19652 7045 182183 7050
rect 19652 6975 20214 7045
rect 20284 6975 182183 7045
rect 19652 6969 182183 6975
rect 182264 6969 182306 7050
rect 533228 6976 533314 6977
rect 540429 6976 540519 6981
rect 533214 6972 540434 6976
rect 182178 6964 182269 6969
rect 180994 6896 181085 6901
rect 533214 6896 533233 6972
rect 533309 6896 540434 6972
rect 540514 6896 540896 6976
rect 180994 6890 180999 6896
rect 19652 6885 180999 6890
rect 19652 6815 20054 6885
rect 20124 6815 180999 6885
rect 181080 6890 181085 6896
rect 533228 6891 533314 6896
rect 540429 6891 540519 6896
rect 181080 6815 181124 6890
rect 535604 6824 535690 6829
rect 535604 6816 535609 6824
rect 19652 6809 181124 6815
rect 535520 6748 535609 6816
rect 535685 6816 535690 6824
rect 540589 6816 540679 6821
rect 535685 6748 540594 6816
rect 178627 6732 178718 6737
rect 535520 6736 540594 6748
rect 540674 6736 540896 6816
rect 178627 6730 178632 6732
rect 19652 6725 178632 6730
rect 19652 6655 19894 6725
rect 19964 6655 178632 6725
rect 19652 6651 178632 6655
rect 178713 6730 178718 6732
rect 540589 6731 540679 6736
rect 178713 6651 178742 6730
rect 540749 6662 540839 6667
rect 540749 6656 540754 6662
rect 19652 6649 178742 6651
rect 178627 6646 178718 6649
rect 536692 6648 540754 6656
rect 177443 6574 177534 6579
rect 536692 6576 536793 6648
rect 177443 6570 177448 6574
rect 19652 6563 177448 6570
rect 19652 6493 19734 6563
rect 19804 6493 177448 6563
rect 177529 6570 177534 6574
rect 536788 6572 536793 6576
rect 536869 6582 540754 6648
rect 540834 6656 540839 6662
rect 540834 6582 540896 6656
rect 536869 6576 540896 6582
rect 536869 6572 536874 6576
rect 177529 6493 177576 6570
rect 536788 6567 536874 6572
rect 539145 6496 539231 6501
rect 565269 6498 565359 6503
rect 565269 6496 565274 6498
rect 19652 6489 177576 6493
rect 19729 6488 19809 6489
rect 177443 6488 177534 6489
rect 539030 6420 539150 6496
rect 539226 6420 565274 6496
rect 539030 6418 565274 6420
rect 565354 6496 565359 6498
rect 565354 6418 565898 6496
rect 539030 6416 565898 6418
rect 539145 6415 539231 6416
rect 565269 6413 565359 6416
rect 175088 6410 175179 6413
rect 18654 6408 175204 6410
rect 18654 6403 175093 6408
rect 18654 6333 19214 6403
rect 19284 6333 175093 6403
rect 18654 6329 175093 6333
rect 19209 6328 19289 6329
rect 175088 6327 175093 6329
rect 175174 6329 175204 6408
rect 565429 6344 565519 6349
rect 565429 6336 565434 6344
rect 175174 6327 175179 6329
rect 175088 6322 175179 6327
rect 540288 6324 565434 6336
rect 540288 6256 540334 6324
rect 19049 6250 19129 6252
rect 173904 6250 173995 6253
rect 18654 6248 174012 6250
rect 18654 6247 173909 6248
rect 18654 6177 19054 6247
rect 19124 6177 173909 6247
rect 18654 6169 173909 6177
rect 173904 6167 173909 6169
rect 173990 6169 174012 6248
rect 540329 6248 540334 6256
rect 540410 6264 565434 6324
rect 565514 6336 565519 6344
rect 565514 6264 565898 6336
rect 540410 6256 565898 6264
rect 540410 6248 540415 6256
rect 540329 6243 540415 6248
rect 565589 6180 565679 6185
rect 542701 6176 542788 6177
rect 565589 6176 565594 6180
rect 542648 6172 565594 6176
rect 173990 6167 173995 6169
rect 173904 6162 173995 6167
rect 171561 6094 171652 6099
rect 542648 6096 542706 6172
rect 171561 6090 171566 6094
rect 18654 6083 171566 6090
rect 18654 6013 18894 6083
rect 18964 6013 171566 6083
rect 171647 6090 171652 6094
rect 542701 6095 542706 6096
rect 542783 6100 565594 6172
rect 565674 6176 565679 6180
rect 565674 6100 565898 6176
rect 542783 6096 565898 6100
rect 542783 6095 542788 6096
rect 565589 6095 565679 6096
rect 542701 6090 542788 6095
rect 171647 6013 171706 6090
rect 543885 6016 543972 6017
rect 565749 6016 565839 6019
rect 18654 6009 171706 6013
rect 543806 6014 565898 6016
rect 543806 6012 565754 6014
rect 18889 6008 18969 6009
rect 171561 6008 171652 6009
rect 543806 5936 543890 6012
rect 543885 5935 543890 5936
rect 543967 5936 565754 6012
rect 543967 5935 543972 5936
rect 170377 5930 170468 5935
rect 543885 5930 543972 5935
rect 565749 5934 565754 5936
rect 565834 5936 565898 6014
rect 584320 5977 585600 6002
rect 565834 5934 565839 5936
rect 18654 5919 170382 5930
rect 18654 5849 18734 5919
rect 18804 5849 170382 5919
rect 170463 5849 170518 5930
rect 565749 5929 565839 5934
rect 584284 5896 585600 5977
rect 584320 5890 585600 5896
rect 546246 5860 546333 5865
rect 546246 5856 546251 5860
rect 18729 5844 18809 5849
rect 170377 5844 170468 5849
rect 546202 5783 546251 5856
rect 546328 5856 546333 5860
rect 566269 5856 566359 5859
rect 546328 5854 566900 5856
rect 546328 5783 566274 5854
rect 546202 5776 566274 5783
rect 566269 5774 566274 5776
rect 566354 5776 566900 5854
rect 566354 5774 566359 5776
rect 167997 5770 168088 5773
rect 17676 5768 168122 5770
rect 566269 5769 566359 5774
rect 17676 5763 168002 5768
rect 17676 5693 18214 5763
rect 18284 5693 168002 5763
rect 17676 5689 168002 5693
rect 18209 5688 18289 5689
rect 167997 5687 168002 5689
rect 168083 5689 168122 5768
rect 547430 5700 547517 5705
rect 547430 5696 547435 5700
rect 168083 5687 168088 5689
rect 167997 5682 168088 5687
rect 547390 5623 547435 5696
rect 547512 5696 547517 5700
rect 566429 5700 566519 5705
rect 566429 5696 566434 5700
rect 547512 5623 566434 5696
rect 547390 5620 566434 5623
rect 566514 5696 566519 5700
rect 566514 5620 566900 5696
rect 547390 5616 566900 5620
rect 566429 5615 566519 5616
rect 18049 5610 18129 5612
rect 166813 5610 166904 5613
rect 17676 5608 166922 5610
rect 17676 5607 166818 5608
rect 17676 5537 18054 5607
rect 18124 5537 166818 5607
rect 17676 5529 166818 5537
rect 166813 5527 166818 5529
rect 166899 5529 166922 5608
rect 566589 5542 566679 5547
rect 566589 5536 566594 5542
rect 166899 5527 166904 5529
rect 166813 5522 166904 5527
rect 549736 5528 566594 5536
rect 549736 5456 549788 5528
rect 549783 5451 549788 5456
rect 549865 5462 566594 5528
rect 566674 5536 566679 5542
rect 566674 5462 566900 5536
rect 549865 5456 566900 5462
rect 549865 5451 549870 5456
rect 164452 5450 164543 5451
rect 17676 5446 164574 5450
rect 549783 5446 549870 5451
rect 17676 5443 164457 5446
rect 17676 5373 17894 5443
rect 17964 5373 164457 5443
rect 17676 5369 164457 5373
rect 17889 5368 17969 5369
rect 164452 5365 164457 5369
rect 164538 5369 164574 5446
rect 566749 5380 566839 5385
rect 550967 5376 551054 5377
rect 566749 5376 566754 5380
rect 550932 5372 566754 5376
rect 164538 5365 164543 5369
rect 164452 5360 164543 5365
rect 163268 5302 163359 5307
rect 163268 5290 163273 5302
rect 17676 5281 163273 5290
rect 17676 5211 17734 5281
rect 17804 5221 163273 5281
rect 163354 5290 163359 5302
rect 550932 5296 550972 5372
rect 550967 5295 550972 5296
rect 551049 5300 566754 5372
rect 566834 5376 566839 5380
rect 566834 5300 566900 5376
rect 551049 5296 566900 5300
rect 551049 5295 551054 5296
rect 566749 5295 566839 5296
rect 550967 5290 551054 5295
rect 163354 5221 163376 5290
rect 17804 5211 163376 5221
rect 553341 5218 553428 5223
rect 553341 5216 553346 5218
rect 17676 5209 163376 5211
rect 17729 5206 17809 5209
rect 553306 5141 553346 5216
rect 553423 5216 553428 5218
rect 567269 5216 567359 5221
rect 553423 5141 567274 5216
rect 553306 5136 567274 5141
rect 567354 5136 567914 5216
rect 567269 5131 567359 5136
rect 16696 5124 161040 5130
rect 16696 5123 160918 5124
rect 16696 5053 17214 5123
rect 17284 5053 160918 5123
rect 16696 5049 160918 5053
rect 17209 5048 17289 5049
rect 160913 5043 160918 5049
rect 160999 5049 161040 5124
rect 567429 5060 567519 5065
rect 567429 5056 567434 5060
rect 160999 5043 161004 5049
rect 160913 5038 161004 5043
rect 554478 5046 567434 5056
rect 554478 4976 554530 5046
rect 16696 4963 159856 4970
rect 554525 4969 554530 4976
rect 554607 4980 567434 5046
rect 567514 5056 567519 5060
rect 567514 4980 567914 5056
rect 554607 4976 567914 4980
rect 554607 4969 554612 4976
rect 567429 4975 567519 4976
rect 554525 4964 554612 4969
rect 16696 4893 17054 4963
rect 17124 4956 159856 4963
rect 17124 4893 159734 4956
rect 16696 4889 159734 4893
rect 17049 4888 17129 4889
rect 159729 4875 159734 4889
rect 159815 4889 159856 4956
rect 567589 4902 567679 4907
rect 556881 4896 556975 4899
rect 567589 4896 567594 4902
rect 556842 4894 567594 4896
rect 159815 4875 159820 4889
rect 159729 4870 159820 4875
rect 800 4708 6370 4820
rect 556842 4816 556886 4894
rect 157355 4810 157446 4811
rect 556881 4810 556886 4816
rect 556970 4822 567594 4894
rect 567674 4896 567679 4902
rect 567674 4822 567914 4896
rect 556970 4816 567914 4822
rect 556970 4810 556975 4816
rect 16696 4806 157472 4810
rect 16696 4799 157360 4806
rect 16696 4729 16894 4799
rect 16964 4729 157360 4799
rect 16889 4724 16969 4729
rect 157355 4725 157360 4729
rect 157441 4729 157472 4806
rect 556881 4805 556975 4810
rect 584320 4797 585600 4820
rect 558065 4736 558159 4739
rect 567749 4736 567839 4737
rect 558000 4734 567914 4736
rect 157441 4725 157446 4729
rect 157355 4720 157446 4725
rect 156171 4652 156262 4657
rect 558000 4656 558070 4734
rect 156171 4650 156176 4652
rect 16696 4637 156176 4650
rect 16696 4569 16734 4637
rect 16729 4567 16734 4569
rect 16804 4571 156176 4637
rect 156257 4650 156262 4652
rect 558065 4650 558070 4656
rect 558154 4732 567914 4734
rect 558154 4656 567754 4732
rect 558154 4650 558159 4656
rect 156257 4571 156286 4650
rect 558065 4645 558159 4650
rect 567749 4652 567754 4656
rect 567834 4656 567914 4732
rect 584284 4730 585600 4797
rect 584320 4708 585600 4730
rect 567834 4652 567839 4656
rect 567749 4647 567839 4652
rect 568269 4576 568359 4579
rect 16804 4569 156286 4571
rect 560372 4574 568890 4576
rect 560372 4571 568274 4574
rect 16804 4567 16809 4569
rect 16729 4562 16809 4567
rect 156171 4566 156262 4569
rect 560372 4501 560425 4571
rect 560495 4501 568274 4571
rect 560372 4496 568274 4501
rect 568269 4494 568274 4496
rect 568354 4496 568890 4574
rect 568354 4494 568359 4496
rect 16209 4490 16289 4494
rect 153803 4490 153894 4493
rect 15650 4489 153928 4490
rect 568269 4489 568359 4494
rect 15650 4419 16214 4489
rect 16284 4488 153928 4489
rect 16284 4419 153808 4488
rect 15650 4409 153808 4419
rect 153803 4407 153808 4409
rect 153889 4409 153928 4488
rect 561528 4411 568890 4416
rect 153889 4407 153894 4409
rect 153803 4402 153894 4407
rect 561528 4341 561625 4411
rect 561695 4408 568890 4411
rect 561695 4341 568434 4408
rect 152619 4334 152710 4339
rect 561528 4336 568434 4341
rect 16049 4330 16129 4332
rect 152619 4330 152624 4334
rect 15650 4327 152624 4330
rect 15650 4257 16054 4327
rect 16124 4257 152624 4327
rect 15650 4253 152624 4257
rect 152705 4330 152710 4334
rect 152705 4253 152742 4330
rect 568429 4328 568434 4336
rect 568514 4336 568890 4408
rect 568514 4328 568519 4336
rect 568429 4323 568519 4328
rect 563975 4262 564061 4267
rect 563975 4256 563980 4262
rect 15650 4249 152742 4253
rect 152619 4248 152710 4249
rect 563934 4186 563980 4256
rect 564056 4256 564061 4262
rect 564056 4250 568890 4256
rect 564056 4186 568594 4250
rect 563934 4176 568594 4186
rect 15889 4170 15969 4172
rect 150277 4170 150368 4175
rect 568589 4170 568594 4176
rect 568674 4176 568890 4250
rect 568674 4170 568679 4176
rect 15650 4167 150282 4170
rect 15650 4097 15894 4167
rect 15964 4097 150282 4167
rect 15650 4089 150282 4097
rect 150363 4089 150394 4170
rect 568589 4165 568679 4170
rect 565159 4102 565245 4107
rect 565159 4096 565164 4102
rect 150277 4084 150368 4089
rect 565118 4026 565164 4096
rect 565240 4096 565245 4102
rect 568749 4096 568839 4097
rect 565240 4092 568890 4096
rect 565240 4026 568754 4092
rect 565118 4016 568754 4026
rect 149093 4010 149184 4013
rect 568749 4012 568754 4016
rect 568834 4016 568890 4092
rect 568834 4012 568839 4016
rect 15650 4008 149228 4010
rect 15650 3999 149098 4008
rect 15650 3929 15734 3999
rect 15804 3929 149098 3999
rect 15729 3924 15809 3929
rect 149093 3927 149098 3929
rect 149179 3929 149228 4008
rect 568749 4007 568839 4012
rect 567522 3941 567610 3946
rect 567522 3936 567527 3941
rect 149179 3927 149184 3929
rect 149093 3922 149184 3927
rect 567468 3863 567527 3936
rect 567605 3936 567610 3941
rect 567605 3924 569916 3936
rect 567605 3863 569274 3924
rect 146719 3852 146810 3857
rect 567468 3856 569274 3863
rect 146719 3850 146724 3852
rect 14680 3841 146724 3850
rect 14680 3771 15214 3841
rect 15284 3771 146724 3841
rect 146805 3850 146810 3852
rect 146805 3771 146822 3850
rect 569269 3844 569274 3856
rect 569354 3856 569916 3924
rect 569354 3844 569359 3856
rect 569269 3839 569359 3844
rect 568706 3776 568794 3778
rect 569429 3776 569519 3777
rect 14680 3769 146822 3771
rect 568664 3773 569916 3776
rect 15209 3766 15289 3769
rect 146719 3766 146810 3769
rect 145535 3694 145626 3699
rect 568664 3696 568711 3773
rect 145535 3690 145540 3694
rect 14680 3685 145540 3690
rect 800 3526 1280 3638
rect 14680 3615 15054 3685
rect 15124 3615 145540 3685
rect 14680 3613 145540 3615
rect 145621 3690 145626 3694
rect 568706 3695 568711 3696
rect 568789 3772 569916 3773
rect 568789 3696 569434 3772
rect 568789 3695 568794 3696
rect 568706 3690 568794 3695
rect 569429 3692 569434 3696
rect 569514 3696 569916 3772
rect 569514 3692 569519 3696
rect 145621 3613 145664 3690
rect 569429 3687 569519 3692
rect 569589 3616 569679 3617
rect 571045 3616 571133 3620
rect 14680 3609 145664 3613
rect 569248 3615 571186 3616
rect 569248 3612 571050 3615
rect 145535 3608 145626 3609
rect 143186 3534 143277 3539
rect 569248 3536 569594 3612
rect 143186 3530 143191 3534
rect 14680 3519 143191 3530
rect 14680 3449 14894 3519
rect 14964 3453 143191 3519
rect 143272 3530 143277 3534
rect 569589 3532 569594 3536
rect 569674 3537 571050 3612
rect 571128 3537 571186 3615
rect 569674 3536 571186 3537
rect 569674 3532 569679 3536
rect 571045 3532 571133 3536
rect 143272 3453 143294 3530
rect 569589 3527 569679 3532
rect 584320 3526 584800 3638
rect 572229 3461 572317 3466
rect 569749 3456 569839 3459
rect 572229 3456 572234 3461
rect 14964 3449 143294 3453
rect 569248 3454 572234 3456
rect 14889 3444 14969 3449
rect 143186 3448 143277 3449
rect 569248 3376 569754 3454
rect 569749 3374 569754 3376
rect 569834 3383 572234 3454
rect 572312 3456 572317 3461
rect 572312 3383 572426 3456
rect 569834 3376 572426 3383
rect 569834 3374 569839 3376
rect 142002 3370 142093 3373
rect 14680 3368 142144 3370
rect 569749 3369 569839 3374
rect 14680 3363 142007 3368
rect 14680 3293 14734 3363
rect 14804 3293 142007 3363
rect 14680 3289 142007 3293
rect 14729 3288 14809 3289
rect 142002 3287 142007 3289
rect 142088 3289 142144 3368
rect 570269 3298 570359 3303
rect 570269 3296 570274 3298
rect 142088 3287 142093 3289
rect 142002 3282 142093 3287
rect 139628 3216 139719 3221
rect 570228 3218 570274 3296
rect 570354 3296 570359 3298
rect 574605 3296 574693 3300
rect 570354 3295 574698 3296
rect 570354 3218 574610 3295
rect 570228 3217 574610 3218
rect 574688 3217 574698 3295
rect 570228 3216 574698 3217
rect 139628 3210 139633 3216
rect 13634 3199 139633 3210
rect 13634 3129 14214 3199
rect 14284 3135 139633 3199
rect 139714 3210 139719 3216
rect 570269 3213 570359 3216
rect 574605 3212 574693 3216
rect 139714 3135 139752 3210
rect 570429 3136 570519 3141
rect 575789 3139 575877 3144
rect 575789 3136 575794 3139
rect 14284 3129 139752 3135
rect 14209 3124 14289 3129
rect 570228 3056 570434 3136
rect 570514 3061 575794 3136
rect 575872 3136 575877 3139
rect 575872 3061 575916 3136
rect 570514 3056 575916 3061
rect 138444 3050 138535 3055
rect 570429 3051 570519 3056
rect 13634 3043 138449 3050
rect 13634 2973 14054 3043
rect 14124 2973 138449 3043
rect 13634 2969 138449 2973
rect 138530 2969 138574 3050
rect 570589 2976 570679 2981
rect 578149 2977 578237 2982
rect 578149 2976 578154 2977
rect 14049 2968 14129 2969
rect 138444 2964 138535 2969
rect 136083 2900 136174 2905
rect 136083 2890 136088 2900
rect 13634 2883 136088 2890
rect 13634 2813 13894 2883
rect 13964 2819 136088 2883
rect 136169 2890 136174 2900
rect 570228 2896 570594 2976
rect 570674 2899 578154 2976
rect 578232 2976 578237 2977
rect 578232 2899 578314 2976
rect 570674 2896 578314 2899
rect 570589 2891 570679 2896
rect 578149 2894 578237 2896
rect 136169 2819 136220 2890
rect 13964 2813 136220 2819
rect 579333 2816 579421 2820
rect 13634 2809 136220 2813
rect 570228 2815 579442 2816
rect 13889 2808 13969 2809
rect 570228 2808 579338 2815
rect 570228 2736 570754 2808
rect 134899 2730 134990 2733
rect 13634 2728 135034 2730
rect 13634 2723 134904 2728
rect 13634 2653 13734 2723
rect 13804 2653 134904 2723
rect 13634 2649 134904 2653
rect 13729 2648 13809 2649
rect 134899 2647 134904 2649
rect 134985 2649 135034 2728
rect 570749 2728 570754 2736
rect 570834 2737 579338 2808
rect 579416 2737 579442 2815
rect 570834 2736 579442 2737
rect 570834 2728 570839 2736
rect 579333 2732 579421 2736
rect 570749 2723 570839 2728
rect 134985 2647 134990 2649
rect 134899 2642 134990 2647
rect 12606 2563 132674 2570
rect 12606 2493 13134 2563
rect 13204 2562 132674 2563
rect 13204 2493 132555 2562
rect 12606 2489 132555 2493
rect 13129 2488 13209 2489
rect 132550 2481 132555 2489
rect 132636 2489 132674 2562
rect 132636 2481 132641 2489
rect 132550 2476 132641 2481
rect 800 2344 1280 2456
rect 12989 2410 13069 2412
rect 131366 2410 131457 2411
rect 12606 2407 131474 2410
rect 12606 2337 12994 2407
rect 13064 2406 131474 2407
rect 13064 2337 131371 2406
rect 12606 2329 131371 2337
rect 131366 2325 131371 2329
rect 131452 2329 131474 2406
rect 584320 2344 584800 2456
rect 131452 2325 131457 2329
rect 131366 2320 131457 2325
rect 128997 2260 129088 2265
rect 12849 2250 12929 2252
rect 128997 2250 129002 2260
rect 12606 2247 129002 2250
rect 12606 2177 12854 2247
rect 12924 2179 129002 2247
rect 129083 2250 129088 2260
rect 129083 2179 129114 2250
rect 12924 2177 129114 2179
rect 12606 2169 129114 2177
rect 127813 2090 127904 2093
rect 12606 2088 127936 2090
rect 12606 2079 127818 2088
rect 12606 2009 12714 2079
rect 12784 2009 127818 2079
rect 12709 2004 12789 2009
rect 127813 2007 127818 2009
rect 127899 2009 127936 2088
rect 127899 2007 127904 2009
rect 127813 2002 127904 2007
<< rmetal3 >>
rect 2884 506420 2996 506532
rect 1988 463198 2100 463310
rect 1780 419976 1892 420088
rect 1810 376754 1922 376866
rect 2154 333532 2266 333644
rect 2144 290310 2256 290422
rect 2464 247288 2576 247400
rect 1558 119666 1678 119778
rect 584048 590572 584160 590684
rect 584088 500850 584200 500962
rect 1310 17710 1430 17822
rect 584000 456428 584112 456540
rect 583888 412006 584000 412118
rect 583886 320362 583998 320474
rect 583996 275940 584108 276052
rect 584076 92372 584180 92484
rect 583772 47714 583894 47826
rect 583772 21256 583898 21368
rect 583488 16528 583600 16640
<< via3 >>
rect 3472 644833 8318 649314
rect 3494 634779 8340 639260
rect 4054 560414 9132 564868
rect 4066 550426 9144 554880
rect 13733 518260 14039 518566
rect 14156 517330 14476 517650
rect 14438 512350 14834 512746
rect 14566 511322 14962 511718
rect 14388 510910 14652 511174
rect 10048 507558 10184 507694
rect 9906 506420 10018 506532
rect 17831 510911 18093 511173
rect 24133 475060 24439 475366
rect 24168 474130 24488 474450
rect 23500 469150 23896 469546
rect 80086 496202 80170 496286
rect 31040 491436 31580 491976
rect 100018 504650 102298 507328
rect 29932 490460 30472 491000
rect 30117 488475 30227 488585
rect 60016 475061 60320 475365
rect 80947 475060 81253 475366
rect 60057 474131 60375 474449
rect 82110 474130 82430 474450
rect 60075 469759 60469 470153
rect 83436 469758 83832 470154
rect 60097 468961 60491 469355
rect 83404 468960 83800 469356
rect 24416 468122 24812 468518
rect 3498 464380 3610 464492
rect 95464 463198 95576 463310
rect 80599 436117 80905 436423
rect 80692 435514 81012 435834
rect 80686 434810 81082 435206
rect 80710 434164 81106 434560
rect 80470 426023 80670 426223
rect 80486 424701 80686 424901
rect 80480 424396 80680 424596
rect 2992 421158 3104 421270
rect 5048 419976 5160 420088
rect 80418 412714 80618 412914
rect 104310 446394 106146 448182
rect 83873 393365 84179 393671
rect 83834 392834 84154 393154
rect 83820 392236 84216 392632
rect 83826 391468 84222 391864
rect 77158 390482 77222 390546
rect 16168 376754 16280 376866
rect 15949 345260 16255 345566
rect 15964 344330 16284 344650
rect 28370 340870 28470 340970
rect 15408 339350 15804 339746
rect 16244 338322 16640 338718
rect 13964 334714 14076 334826
rect 14124 333532 14236 333644
rect 15156 307378 15420 307642
rect 13889 302060 14195 302366
rect 14130 301130 14450 301450
rect 13166 296150 13562 296546
rect 69415 376755 69525 376865
rect 72878 376754 72990 376866
rect 71906 352064 72018 352176
rect 44239 334472 44745 334978
rect 44253 333578 44735 334060
rect 16765 307379 17027 307641
rect 32495 295645 32673 295823
rect 13890 295122 14286 295518
rect 31883 294739 32061 294917
rect 66377 283675 67967 285265
rect 14880 281572 15184 281876
rect 66223 281571 66529 281877
rect 15615 280815 15933 281133
rect 66290 280814 66610 281134
rect 77941 389853 78075 389987
rect 77158 279466 77222 279530
rect 78789 388939 79199 389349
rect 77158 278282 77222 278346
rect 66317 276361 67907 277951
rect 32500 274181 32680 274361
rect 31882 273881 32062 274061
rect 14879 259060 15185 259366
rect 15614 258130 15934 258450
rect 15582 253150 15978 253546
rect 14736 252122 15132 252518
rect 11476 247288 11588 247400
rect 4310 215890 9440 220396
rect 13573 247289 13683 247399
rect 69747 223542 70409 224204
rect 69873 222730 70535 223392
rect 4284 205852 9414 210358
rect 3756 173829 8602 178310
rect 3676 163839 8522 168320
rect 79990 388105 80235 388350
rect 78004 132506 79115 133617
rect 22349 131638 22655 131944
rect 78265 131168 78643 131546
rect 23322 130708 23642 131028
rect 23176 125728 23572 126124
rect 23194 124700 23590 125096
rect 78253 128787 78631 129165
rect 47794 126745 48905 127856
rect 77898 119666 78010 119778
rect 116072 345626 118072 347766
rect 130013 612731 131571 614289
rect 136986 639691 140674 644370
rect 137993 597505 139391 598903
rect 129074 589599 132598 595069
rect 127105 496203 127187 496285
rect 122182 284192 124562 286830
rect 130223 563816 131253 564299
rect 131253 563816 131421 564299
rect 130223 563101 131421 563816
rect 130494 520554 130798 520558
rect 130494 520258 130498 520554
rect 130498 520258 130794 520554
rect 130794 520258 130798 520554
rect 130494 520254 130798 520258
rect 130371 490461 130909 490999
rect 130662 481298 130966 481602
rect 129018 475062 132644 478334
rect 129018 473816 130159 475062
rect 130159 473816 131405 475062
rect 131405 473816 132644 475062
rect 129018 472030 132644 473816
rect 130729 463199 130839 463309
rect 130708 436118 131012 436422
rect 130461 424397 130659 424595
rect 130591 412715 130789 412913
rect 130804 393366 131108 393670
rect 128918 379827 132762 380144
rect 128962 376582 132722 377026
rect 128893 363838 132628 364692
rect 130472 355822 130776 356126
rect 130656 334473 131160 334977
rect 128934 310102 132738 310649
rect 130624 302061 130928 302365
rect 130802 279254 131106 279558
rect 29441 88438 29747 88744
rect 29646 87508 29966 87828
rect 29596 82528 29992 82924
rect 29604 81500 30000 81896
rect 120566 80948 120962 81344
rect 42786 58139 44174 59527
rect 24125 45238 24431 45544
rect 24086 44308 24406 44628
rect 23432 39328 23828 39724
rect 23402 38300 23798 38696
rect 120567 40933 120961 41327
rect 130162 234296 130822 234956
rect 129023 168834 132621 173511
rect 130688 136524 130992 136828
rect 130506 131169 130882 131545
rect 130809 119667 130919 119777
rect 129090 115062 132624 119218
rect 129090 113816 130007 115062
rect 130007 113816 131253 115062
rect 131253 113816 132624 115062
rect 129090 112664 132624 113816
rect 130670 88439 130974 88743
rect 130143 45059 131729 46645
rect 130662 43772 130966 44076
rect 138121 572158 139319 573356
rect 138459 519501 138777 519505
rect 138459 519191 138463 519501
rect 138463 519191 138773 519501
rect 138773 519191 138777 519501
rect 138459 519187 138777 519191
rect 138631 491437 139169 491975
rect 138317 480181 138635 480499
rect 138711 435515 139029 435833
rect 138589 424702 138787 424900
rect 138495 404349 138813 404667
rect 137099 391475 140611 401010
rect 136999 378850 140729 379269
rect 136912 361328 140668 362468
rect 138801 354675 139119 354993
rect 138718 333579 139198 334059
rect 136918 309106 140746 309624
rect 138483 301131 138801 301449
rect 138369 278233 138687 278551
rect 138658 233036 139318 233696
rect 146008 143960 148318 146268
rect 138813 135715 139131 136033
rect 138734 128788 139110 129164
rect 138953 87509 139271 87827
rect 511510 693868 516020 698944
rect 521554 693856 526064 698932
rect 422844 604042 425668 606998
rect 426592 428204 428498 430286
rect 427136 284006 430734 287604
rect 444374 635697 448011 640383
rect 445990 598724 446366 599100
rect 445999 591873 446317 592191
rect 446115 516171 446433 516489
rect 445899 511073 446217 511391
rect 445837 495187 446155 495191
rect 445837 494877 445841 495187
rect 445841 494877 446151 495187
rect 446151 494877 446155 495187
rect 445837 494873 446155 494877
rect 445803 492239 446025 492461
rect 445789 481969 446107 482287
rect 573828 640732 578952 645170
rect 573842 630762 578966 635200
rect 493997 604985 495991 606979
rect 453800 597850 454176 598226
rect 509749 603455 510127 603833
rect 509797 602495 510175 602873
rect 498783 595339 500777 597333
rect 454030 593103 454334 593107
rect 454030 592807 454034 593103
rect 454034 592807 454330 593103
rect 454330 592807 454334 593103
rect 454030 592803 454334 592807
rect 564589 592802 564895 593108
rect 564650 591872 564970 592192
rect 584048 599516 584160 599628
rect 564510 586892 564906 587288
rect 564428 585864 564824 586260
rect 575644 551600 580768 556038
rect 575630 541566 580754 546004
rect 523953 528823 524507 529377
rect 524038 528018 524358 528338
rect 524166 527410 524486 527730
rect 524150 526285 524711 526846
rect 454037 515279 454355 515597
rect 453982 512003 454286 512307
rect 561367 512002 561673 512308
rect 561436 511072 561756 511392
rect 561334 506092 561730 506488
rect 561382 505064 561778 505460
rect 583162 504652 583426 504916
rect 582282 503772 582442 503932
rect 559848 502678 559960 502790
rect 453846 495803 454150 496107
rect 454027 489805 454225 490003
rect 454076 483336 454380 483340
rect 454076 483040 454080 483336
rect 454080 483040 454376 483336
rect 454376 483040 454380 483336
rect 454076 483036 454380 483040
rect 451714 390482 451778 390546
rect 451236 389852 451372 389988
rect 450424 388938 450836 389350
rect 442634 386487 443287 387140
rect 439833 385293 439963 385423
rect 439337 383041 439555 383259
rect 438563 382294 438742 382473
rect 441444 383887 442145 384588
rect 449325 387917 449759 388351
rect 561171 495802 561477 496108
rect 583163 496017 583425 496279
rect 561240 494872 561560 495192
rect 543806 492238 544030 492462
rect 542206 489804 542406 490004
rect 528282 488997 528711 489426
rect 560790 489892 561186 490288
rect 560722 488864 561118 489260
rect 561780 488448 562108 488776
rect 583194 488452 583458 488716
rect 581531 485911 581617 485997
rect 487304 480314 487700 480710
rect 486350 479056 486746 479452
rect 556419 479202 556725 479508
rect 562984 479203 563288 479507
rect 556614 478272 556934 478592
rect 563127 478273 563445 478591
rect 537940 476978 538369 477407
rect 487305 473293 487699 473687
rect 486351 472265 486745 472659
rect 483617 470965 483727 471075
rect 570859 479202 571165 479508
rect 583753 479269 583863 479379
rect 570852 478272 571172 478592
rect 570704 473292 571100 473688
rect 570720 472264 571116 472660
rect 582282 471852 582546 472116
rect 505921 390191 506251 390521
rect 446017 316873 446335 317191
rect 444618 301612 447812 310980
rect 446021 277673 446339 277991
rect 445726 244170 446099 244543
rect 431353 163637 434495 167041
rect 444303 179958 448071 180774
rect 452461 373109 455428 376076
rect 545330 373108 548299 376077
rect 453990 317803 454294 318107
rect 452458 295062 455712 299098
rect 452458 293816 453707 295062
rect 453707 293816 454953 295062
rect 454953 293816 455712 295062
rect 452458 292718 455712 293816
rect 453710 278603 454014 278907
rect 477612 283320 477920 283628
rect 563802 261374 563878 261450
rect 563738 256896 563814 256972
rect 563752 255360 563828 255436
rect 453947 245207 454265 245525
rect 452333 187251 455990 191899
rect 452276 176624 456058 177478
rect 444290 91356 448055 92247
rect 446267 74534 446558 74825
rect 159964 63802 162104 66158
rect 436136 63691 439734 67289
rect 137772 58139 139160 59527
rect 452241 88492 456105 89388
rect 453466 73571 453843 73948
rect 477769 252435 478308 252974
rect 476829 247477 477147 247795
rect 138597 42905 138915 43223
rect 137083 31547 140503 40865
rect 3562 17264 4344 18157
rect 124736 17233 125692 18189
rect 462586 245206 462906 245526
rect 462667 244169 463042 244544
rect 580504 470964 580616 471076
rect 583752 456946 583864 457058
rect 583195 451647 583457 451909
rect 583228 412006 583340 412118
rect 581532 410854 581616 410938
rect 582283 407261 582545 407523
rect 577998 346082 580967 349051
rect 571149 317802 571455 318108
rect 582955 319193 583029 319267
rect 571168 316872 571488 317192
rect 582511 315523 582773 315785
rect 571054 311892 571450 312288
rect 571068 310864 571464 311260
rect 582510 310452 582774 310716
rect 531657 185114 531892 185349
rect 532235 185174 532470 185409
rect 532835 185322 533054 185541
rect 571467 278602 571773 278908
rect 571458 277672 571778 277992
rect 582687 276053 582761 276127
rect 583490 276052 583566 276128
rect 583253 274783 583327 274857
rect 571326 272692 571722 273088
rect 571282 271664 571678 272060
rect 533414 179406 533635 179627
rect 532234 161712 532471 161949
rect 510864 151142 511157 151435
rect 511041 150369 511420 150748
rect 510809 149297 511483 149971
rect 511010 148158 511630 148778
rect 551029 148159 551647 148777
rect 532834 81185 533055 81406
rect 574934 236252 580058 240690
rect 574962 226222 580086 230660
rect 574896 192412 580020 196850
rect 574908 182368 580032 186806
rect 575156 147818 580280 152256
rect 575102 137756 580226 142194
rect 560528 93493 560747 93712
rect 531656 63534 531893 63771
rect 527286 54956 527579 55249
rect 527333 54353 527712 54732
rect 527695 53335 528369 54009
rect 527852 52256 528472 52876
rect 552581 52257 553199 52875
rect 532272 48896 532384 49008
rect 532878 22438 532990 22550
rect 459576 17233 460532 18189
rect 531698 17710 531810 17822
<< metal4 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 511354 698944 526180 699076
rect 511354 693868 511510 698944
rect 516020 698932 526180 698944
rect 516020 693868 516456 698932
rect 511354 693856 516456 693868
rect 520966 693856 521554 698932
rect 526064 693856 526180 698932
rect 511354 693672 526180 693856
rect 3308 649314 8544 649486
rect 3308 644833 3472 649314
rect 8318 644833 8544 649314
rect 3308 644534 8544 644833
rect 573700 645170 579138 645386
rect 3308 644370 141468 644534
rect 3308 639691 136986 644370
rect 140674 639691 141468 644370
rect 573700 640732 573828 645170
rect 578952 640732 579138 645170
rect 573700 640538 579138 640732
rect 3308 639534 141468 639691
rect 443754 640383 579138 640538
rect 3308 639260 8544 639534
rect 3308 634779 3494 639260
rect 8340 634779 8544 639260
rect 443754 635697 444374 640383
rect 448011 635697 579138 640383
rect 443754 635538 579138 635697
rect 3308 634618 8544 634779
rect 573700 635200 579138 635538
rect 573700 630762 573842 635200
rect 578966 630762 579138 635200
rect 573700 630566 579138 630762
rect 93380 614289 131572 614290
rect 93380 612731 130013 614289
rect 131571 612731 131572 614289
rect 93380 612730 131572 612731
rect 93380 601578 94940 612730
rect 71902 600018 94940 601578
rect 98259 601186 169654 610368
rect 417050 606998 478782 610324
rect 417050 604042 422844 606998
rect 425668 606979 478782 606998
rect 493996 606979 495992 606980
rect 425668 604985 493997 606979
rect 495991 604985 495992 606979
rect 425668 604042 478782 604985
rect 493996 604984 495992 604985
rect 72108 598134 107279 599819
rect 118297 597983 119982 601186
rect 72108 596298 119982 597983
rect 124082 598903 139392 598904
rect 124082 597505 137993 598903
rect 139391 597505 139392 598903
rect 124082 597504 139392 597505
rect 124082 596096 125482 597504
rect 71718 594696 125482 596096
rect 128823 595069 132844 595370
rect 128823 593559 129074 595069
rect 98259 592599 129074 593559
rect 73684 588596 119472 590281
rect 128823 589599 129074 592599
rect 132598 589599 132844 595069
rect 128823 589258 132844 589599
rect 73684 586760 107507 588445
rect 117787 587297 119472 588596
rect 143715 587297 145836 601186
rect 417050 601142 478782 604042
rect 509748 603833 510128 603834
rect 495753 603455 509749 603833
rect 510127 603455 510128 603833
rect 495753 599101 496131 603455
rect 509748 603454 510128 603455
rect 509796 602873 510176 602874
rect 445989 599100 496131 599101
rect 445989 598724 445990 599100
rect 446366 598724 496131 599100
rect 445989 598723 496131 598724
rect 496845 602495 509797 602873
rect 510175 602718 510176 602873
rect 510175 602606 511130 602718
rect 510175 602495 510176 602606
rect 496845 598227 497223 602495
rect 509796 602494 510176 602495
rect 511018 599628 511130 602606
rect 584047 599628 584161 599629
rect 511018 599516 584048 599628
rect 584160 599516 584161 599628
rect 584047 599515 584161 599516
rect 453799 598226 497223 598227
rect 453799 597850 453800 598226
rect 454176 597850 497223 598226
rect 453799 597849 497223 597850
rect 498782 597333 500778 597334
rect 471323 595339 498783 597333
rect 500777 595339 500778 597333
rect 498782 595338 500778 595339
rect 564588 593108 564896 593109
rect 454029 593107 564589 593108
rect 454029 592803 454030 593107
rect 454334 592803 564589 593107
rect 454029 592802 564589 592803
rect 564895 592802 564896 593108
rect 564588 592801 564896 592802
rect 564649 592192 564971 592193
rect 445998 592191 564650 592192
rect 445998 591873 445999 592191
rect 446317 591873 564650 592191
rect 445998 591872 564650 591873
rect 564970 591872 564971 592192
rect 564649 591871 564971 591872
rect 117787 585612 145836 587297
rect 564509 587288 564907 587289
rect 430778 586892 564510 587288
rect 564906 586892 564907 587288
rect 564509 586891 564907 586892
rect 564427 586260 564825 586261
rect 469808 585864 564428 586260
rect 564824 585864 564825 586260
rect 564427 585863 564825 585864
rect 73684 579654 107787 581339
rect 144031 579503 145836 585612
rect 73684 577818 145836 579503
rect 73888 573356 139320 573357
rect 73888 572158 138121 573356
rect 139319 572158 139320 573356
rect 73888 572157 139320 572158
rect 144151 571794 145836 577818
rect 73888 570109 145836 571794
rect 73888 568273 108171 569958
rect 73888 566785 125938 567985
rect 3906 564868 9344 565044
rect 3906 560414 4054 564868
rect 9132 560414 9344 564868
rect 124738 564300 125938 566785
rect 124738 564299 131422 564300
rect 124738 563101 130223 564299
rect 131421 563101 131422 564299
rect 124738 563100 131422 563101
rect 3906 560048 9344 560414
rect 3906 555362 4066 560048
rect 9170 555362 9344 560048
rect 3906 554880 9344 555362
rect 3906 550426 4066 554880
rect 9144 550426 9344 554880
rect 3906 550224 9344 550426
rect 466125 560021 473749 560331
rect 466125 553646 466599 560021
rect 473439 553646 473749 560021
rect 466125 530621 473749 553646
rect 575502 556038 580940 556170
rect 575502 551600 575644 556038
rect 580768 551600 580940 556038
rect 575502 550970 580940 551600
rect 575502 546532 575622 550970
rect 580746 546532 580940 550970
rect 575502 546004 580940 546532
rect 575502 541566 575630 546004
rect 580754 541566 580940 546004
rect 575502 541350 580940 541566
rect 466125 523885 466547 530621
rect 473413 529377 473749 530621
rect 523952 529377 524508 529378
rect 473413 528823 523953 529377
rect 524507 528823 524508 529377
rect 473413 523885 473749 528823
rect 523952 528822 524508 528823
rect 524037 528338 524359 528339
rect 466125 523522 473749 523885
rect 486192 528018 524038 528338
rect 524358 528018 524359 528338
rect 27731 520558 130799 520559
rect 27731 520254 130494 520558
rect 130798 520254 130799 520558
rect 27731 520253 130799 520254
rect 13732 518566 14040 518567
rect 27731 518566 28037 520253
rect 13732 518260 13733 518566
rect 14039 518260 28037 518566
rect 28648 519505 138778 519506
rect 28648 519187 138459 519505
rect 138777 519187 138778 519505
rect 28648 519186 138778 519187
rect 13732 518259 14040 518260
rect 14155 517650 14477 517651
rect 28648 517650 28968 519186
rect 14155 517330 14156 517650
rect 14476 517330 28968 517650
rect 29672 518376 154256 518772
rect 14155 517329 14477 517330
rect 14437 512746 14835 512747
rect 29672 512746 30068 518376
rect 14437 512350 14438 512746
rect 14834 512350 30068 512746
rect 30630 517542 109858 517938
rect 14437 512349 14835 512350
rect 14565 511718 14963 511719
rect 30630 511718 31026 517542
rect 46652 516805 93040 517146
rect 46652 516258 46993 516805
rect 50527 516004 87782 516401
rect 14565 511322 14566 511718
rect 14962 511322 31026 511718
rect 14565 511321 14963 511322
rect 14387 511174 14653 511175
rect 14387 510910 14388 511174
rect 14652 511173 18094 511174
rect 14652 510911 17831 511173
rect 18093 510911 18094 511173
rect 14652 510910 18094 510911
rect 14387 510909 14653 510910
rect 10047 507694 10185 507695
rect 10047 507558 10048 507694
rect 10184 507558 27382 507694
rect 10047 507557 10185 507558
rect 9905 506532 10019 506533
rect 9905 506420 9906 506532
rect 10018 506420 24864 506532
rect 9905 506419 10019 506420
rect 24752 488586 24864 506420
rect 27246 490238 27382 507558
rect 87385 498127 87782 516004
rect 92699 510368 93040 516805
rect 486192 516490 486512 528018
rect 524037 528017 524359 528018
rect 524165 527730 524487 527731
rect 446114 516489 486512 516490
rect 446114 516171 446115 516489
rect 446433 516171 486512 516489
rect 446114 516170 486512 516171
rect 486772 527410 524166 527730
rect 524486 527410 524487 527730
rect 486772 515598 487092 527410
rect 524165 527409 524487 527410
rect 524149 526846 524712 526847
rect 454036 515597 487092 515598
rect 454036 515279 454037 515597
rect 454355 515279 487092 515597
rect 454036 515278 487092 515279
rect 489160 526285 524150 526846
rect 524711 526285 524712 526846
rect 417050 513709 440192 514324
rect 489160 513709 489721 526285
rect 524149 526284 524712 526285
rect 417050 513148 489721 513709
rect 91502 507328 169654 510368
rect 91502 504650 100018 507328
rect 102298 504650 169654 507328
rect 417050 505142 440192 513148
rect 453950 512308 454338 512346
rect 561366 512308 561674 512309
rect 453950 512307 561367 512308
rect 453950 512003 453982 512307
rect 454286 512003 561367 512307
rect 453950 512002 561367 512003
rect 561673 512002 561674 512308
rect 453950 511966 454338 512002
rect 561366 512001 561674 512002
rect 561435 511392 561757 511393
rect 445898 511391 561436 511392
rect 445898 511073 445899 511391
rect 446217 511073 561436 511391
rect 445898 511072 561436 511073
rect 561756 511072 561757 511392
rect 561435 511071 561757 511072
rect 561333 506488 561731 506489
rect 443122 506092 561334 506488
rect 561730 506092 561731 506488
rect 91502 501186 169654 504650
rect 443122 503768 443518 506092
rect 561333 506091 561731 506092
rect 561381 505460 561779 505461
rect 469780 505064 561382 505460
rect 561778 505064 561779 505460
rect 561381 505063 561779 505064
rect 583161 504916 583427 504917
rect 583161 504652 583162 504916
rect 583426 504652 583427 504916
rect 583161 504651 583427 504652
rect 582281 503932 582443 503933
rect 582281 503772 582282 503932
rect 582442 503772 582443 503932
rect 582281 503771 582443 503772
rect 430838 503372 443518 503768
rect 559847 502790 559961 502791
rect 559847 502678 559848 502790
rect 559960 502678 559961 502790
rect 559847 502677 559961 502678
rect 87385 497730 109971 498127
rect 80085 496286 80171 496287
rect 80085 496202 80086 496286
rect 80170 496285 127188 496286
rect 80170 496203 127105 496285
rect 127187 496203 127188 496285
rect 80170 496202 127188 496203
rect 80085 496201 80171 496202
rect 559848 496108 559960 502677
rect 561170 496108 561478 496109
rect 453845 496107 561171 496108
rect 453845 495803 453846 496107
rect 454150 495803 561171 496107
rect 453845 495802 561171 495803
rect 561477 495802 561478 496108
rect 561170 495801 561478 495802
rect 561239 495192 561561 495193
rect 445836 495191 561240 495192
rect 445836 494873 445837 495191
rect 446155 494873 561240 495191
rect 445836 494872 561240 494873
rect 561560 494872 561561 495192
rect 561239 494871 561561 494872
rect 543805 492462 544031 492463
rect 445802 492461 543806 492462
rect 445802 492239 445803 492461
rect 446025 492239 543806 492461
rect 445802 492238 543806 492239
rect 544030 492238 544031 492462
rect 543805 492237 544031 492238
rect 31039 491976 31581 491977
rect 31039 491436 31040 491976
rect 31580 491975 139170 491976
rect 31580 491437 138631 491975
rect 139169 491437 139170 491975
rect 31580 491436 139170 491437
rect 31039 491435 31581 491436
rect 430344 491342 553364 491738
rect 29931 491000 30473 491001
rect 29931 490460 29932 491000
rect 30472 490999 130994 491000
rect 30472 490461 130371 490999
rect 130909 490461 130994 490999
rect 30472 490460 130994 490461
rect 29931 490459 30473 490460
rect 470194 490244 552214 490640
rect 27246 490102 72602 490238
rect 24752 488585 30250 488586
rect 24752 488475 30117 488585
rect 30227 488475 30250 488585
rect 24752 488474 30250 488475
rect 24132 475366 24440 475367
rect 24132 475060 24133 475366
rect 24439 475365 60321 475366
rect 24439 475061 60016 475365
rect 60320 475061 60321 475365
rect 24439 475060 60321 475061
rect 24132 475059 24440 475060
rect 24167 474450 24489 474451
rect 24167 474130 24168 474450
rect 24488 474449 60376 474450
rect 24488 474131 60057 474449
rect 60375 474131 60376 474449
rect 24488 474130 60376 474131
rect 24167 474129 24489 474130
rect 23500 470153 60470 470154
rect 23500 469759 60075 470153
rect 60469 469759 60470 470153
rect 23500 469758 60470 469759
rect 23500 469547 23896 469758
rect 23499 469546 23897 469547
rect 23499 469150 23500 469546
rect 23896 469150 23897 469546
rect 23499 469149 23897 469150
rect 24416 469355 60492 469356
rect 24416 468961 60097 469355
rect 60491 468961 60492 469355
rect 24416 468960 60492 468961
rect 24416 468519 24812 468960
rect 24415 468518 24813 468519
rect 24415 468122 24416 468518
rect 24812 468122 24813 468518
rect 24415 468121 24813 468122
rect 3497 464492 3611 464493
rect 3497 464380 3498 464492
rect 3610 464380 72038 464492
rect 3497 464379 3611 464380
rect 2991 421270 3105 421271
rect 2991 421158 2992 421270
rect 3104 421158 31168 421270
rect 2991 421157 3105 421158
rect 5047 420088 5161 420089
rect 5047 419976 5048 420088
rect 5160 419976 30194 420088
rect 5047 419975 5161 419976
rect 30082 403922 30194 419976
rect 31056 404788 31168 421158
rect 31056 404676 71446 404788
rect 30082 403810 66926 403922
rect 16167 376866 16281 376867
rect 66814 376866 66926 403810
rect 71334 384588 71446 404676
rect 71926 385423 72038 464380
rect 72466 387140 72602 490102
rect 542205 490004 542407 490005
rect 454026 490003 542206 490004
rect 454026 489805 454027 490003
rect 454225 489805 542206 490003
rect 454026 489804 542206 489805
rect 542406 489804 542407 490004
rect 542205 489803 542407 489804
rect 528281 489426 528712 489427
rect 469600 488997 469678 489426
rect 470107 488997 528282 489426
rect 528711 488997 528712 489426
rect 528281 488996 528712 488997
rect 551818 489260 552214 490244
rect 552968 490288 553364 491342
rect 560789 490288 561187 490289
rect 552968 489892 560790 490288
rect 561186 489892 561187 490288
rect 560789 489891 561187 489892
rect 560721 489260 561119 489261
rect 551818 488864 560722 489260
rect 561118 488864 561119 489260
rect 560721 488863 561119 488864
rect 561779 488776 562109 488777
rect 561779 488448 561780 488776
rect 562108 488448 562109 488776
rect 454075 483340 490027 483341
rect 454075 483036 454076 483340
rect 454380 483036 490027 483340
rect 454075 483035 490027 483036
rect 445788 482287 489176 482288
rect 445788 481969 445789 482287
rect 446107 481969 489176 482287
rect 445788 481968 489176 481969
rect 80947 481602 130967 481603
rect 80947 481298 130662 481602
rect 130966 481298 130967 481602
rect 80947 481297 130967 481298
rect 80947 475367 81253 481297
rect 487303 480710 487701 480711
rect 82110 480499 138636 480500
rect 82110 480181 138317 480499
rect 138635 480181 138636 480499
rect 430596 480314 487304 480710
rect 487700 480314 487701 480710
rect 487303 480313 487701 480314
rect 82110 480180 138636 480181
rect 80946 475366 81254 475367
rect 80946 475060 80947 475366
rect 81253 475060 81254 475366
rect 80946 475059 81254 475060
rect 82110 474451 82430 480180
rect 83436 479222 154442 479618
rect 486349 479452 486747 479453
rect 82109 474450 82431 474451
rect 82109 474130 82110 474450
rect 82430 474130 82431 474450
rect 82109 474129 82431 474130
rect 83436 470155 83832 479222
rect 470690 479056 486350 479452
rect 486746 479056 486747 479452
rect 486349 479055 486747 479056
rect 488856 478592 489176 481968
rect 489721 479508 490027 483035
rect 556418 479508 556726 479509
rect 489721 479202 556419 479508
rect 556725 479202 556726 479508
rect 556418 479201 556726 479202
rect 556613 478592 556935 478593
rect 128648 478334 280759 478540
rect 88986 475380 114425 475493
rect 88986 470556 106611 475380
rect 87180 470309 106611 470556
rect 113894 470309 114425 475380
rect 128648 472030 129018 478334
rect 132644 478254 280759 478334
rect 488856 478272 556614 478592
rect 556934 478272 556935 478592
rect 556613 478271 556935 478272
rect 132644 472070 273502 478254
rect 280420 472070 280759 478254
rect 537939 477407 538370 477408
rect 132644 472030 280759 472070
rect 128648 471802 280759 472030
rect 477920 476978 537940 477407
rect 538369 476978 538370 477407
rect 87180 470219 114425 470309
rect 87180 470160 89804 470219
rect 83435 470154 83833 470155
rect 83435 469758 83436 470154
rect 83832 469758 83833 470154
rect 83435 469757 83833 469758
rect 83403 469356 83801 469357
rect 87180 469356 87576 470160
rect 83403 468960 83404 469356
rect 83800 468960 87576 469356
rect 83403 468959 83801 468960
rect 95463 463310 95577 463311
rect 95463 463198 95464 463310
rect 95576 463309 130840 463310
rect 95576 463199 130729 463309
rect 130839 463199 130840 463309
rect 95576 463198 130840 463199
rect 95463 463197 95577 463198
rect 150797 462824 158032 462940
rect 150797 462028 150899 462824
rect 88986 461395 150899 462028
rect 157916 462028 158032 462824
rect 157916 461395 158180 462028
rect 88986 461302 158180 461395
rect 150797 461301 158032 461302
rect 106510 455757 114021 455761
rect 88986 455661 114021 455757
rect 88986 455031 106619 455661
rect 106510 454319 106619 455031
rect 113903 454319 114021 455661
rect 106510 454196 114021 454319
rect 88986 448182 169654 452168
rect 88986 446394 104310 448182
rect 106146 446394 169654 448182
rect 88986 442986 169654 446394
rect 106528 441575 114020 441685
rect 106528 440841 106630 441575
rect 88986 440408 106630 440841
rect 113902 440841 114020 441575
rect 113902 440408 114120 440841
rect 88986 440326 114120 440408
rect 150780 440395 158029 440524
rect 106528 440321 114020 440326
rect 150780 439439 150941 440395
rect 88986 439040 150941 439439
rect 157881 439040 158029 440395
rect 88986 438906 158029 439040
rect 88986 438904 157979 438906
rect 80598 436423 80906 436424
rect 80598 436117 80599 436423
rect 80905 436422 131013 436423
rect 80905 436118 130708 436422
rect 131012 436118 131013 436422
rect 80905 436117 131013 436118
rect 80598 436116 80906 436117
rect 80691 435834 81013 435835
rect 80691 435514 80692 435834
rect 81012 435833 139030 435834
rect 81012 435515 138711 435833
rect 139029 435515 139030 435833
rect 81012 435514 139030 435515
rect 80691 435513 81013 435514
rect 80685 435206 81083 435207
rect 80685 434810 80686 435206
rect 81082 434810 153732 435206
rect 80685 434809 81083 434810
rect 80709 434560 81107 434561
rect 80709 434164 80710 434560
rect 81106 434164 109890 434560
rect 80709 434163 81107 434164
rect 80469 426223 80671 426224
rect 163014 426223 163214 442986
rect 80469 426023 80470 426223
rect 80670 426023 163214 426223
rect 417050 430286 440192 434324
rect 417050 428204 426592 430286
rect 428498 429993 440192 430286
rect 477920 429993 478349 476978
rect 537939 476977 538370 476978
rect 561779 476233 562109 488448
rect 581530 485997 581618 485998
rect 581530 485911 581531 485997
rect 581617 485911 581618 485997
rect 581530 485910 581618 485911
rect 570858 479508 571166 479509
rect 562983 479507 570859 479508
rect 562983 479203 562984 479507
rect 563288 479203 570859 479507
rect 562983 479202 570859 479203
rect 571165 479202 571166 479508
rect 570858 479201 571166 479202
rect 570851 478592 571173 478593
rect 563126 478591 570852 478592
rect 563126 478273 563127 478591
rect 563445 478273 570852 478591
rect 563126 478272 570852 478273
rect 571172 478272 571173 478592
rect 570851 478271 571173 478272
rect 428498 429564 478349 429993
rect 480469 475903 562109 476233
rect 428498 428204 440192 429564
rect 80469 426022 80671 426023
rect 417050 425142 440192 428204
rect 80485 424901 80687 424902
rect 80485 424701 80486 424901
rect 80686 424900 138788 424901
rect 80686 424702 138589 424900
rect 138787 424702 138788 424900
rect 80686 424701 138788 424702
rect 80485 424700 80687 424701
rect 80479 424596 80681 424597
rect 80479 424396 80480 424596
rect 80680 424595 130660 424596
rect 80680 424397 130461 424595
rect 130659 424397 130660 424595
rect 80680 424396 130660 424397
rect 80479 424395 80681 424396
rect 80417 412914 80619 412915
rect 80417 412714 80418 412914
rect 80618 412913 130790 412914
rect 80618 412715 130591 412913
rect 130789 412715 130790 412913
rect 80618 412714 130790 412715
rect 80417 412713 80619 412714
rect 133778 404667 138814 404668
rect 133778 404349 138495 404667
rect 138813 404349 138814 404667
rect 133778 404348 138814 404349
rect 83872 393671 84180 393672
rect 83872 393365 83873 393671
rect 84179 393670 131109 393671
rect 84179 393366 130804 393670
rect 131108 393366 131109 393670
rect 84179 393365 131109 393366
rect 83872 393364 84180 393365
rect 83833 393154 84155 393155
rect 133778 393154 134098 404348
rect 83833 392834 83834 393154
rect 84154 392834 134098 393154
rect 134706 402698 154300 403094
rect 83833 392833 84155 392834
rect 83819 392632 84217 392633
rect 134706 392632 135102 402698
rect 83819 392236 83820 392632
rect 84216 392236 135102 392632
rect 136611 401010 167867 401173
rect 83819 392235 84217 392236
rect 83825 391864 84223 391865
rect 83825 391468 83826 391864
rect 84222 391468 109920 391864
rect 136611 391475 137099 401010
rect 140611 400684 167867 401010
rect 140611 391614 163821 400684
rect 167356 391614 167867 400684
rect 140611 391475 167867 391614
rect 83825 391467 84223 391468
rect 136611 391172 167867 391475
rect 77157 390546 77223 390547
rect 77157 390482 77158 390546
rect 77222 390544 77223 390546
rect 451713 390546 451779 390547
rect 451713 390544 451714 390546
rect 77222 390484 451714 390544
rect 77222 390482 77223 390484
rect 77157 390481 77223 390482
rect 451713 390482 451714 390484
rect 451778 390482 451779 390546
rect 451713 390481 451779 390482
rect 480469 390521 480799 475903
rect 570703 473688 571101 473689
rect 487304 473687 570704 473688
rect 487304 473293 487305 473687
rect 487699 473293 570704 473687
rect 487304 473292 570704 473293
rect 571100 473292 571101 473688
rect 570703 473291 571101 473292
rect 570719 472660 571117 472661
rect 486350 472659 570720 472660
rect 486350 472265 486351 472659
rect 486745 472265 570720 472659
rect 486350 472264 570720 472265
rect 571116 472264 571117 472660
rect 570719 472263 571117 472264
rect 580503 471076 580617 471077
rect 483616 471075 580504 471076
rect 483616 470965 483617 471075
rect 483727 470965 580504 471075
rect 483616 470964 580504 470965
rect 580616 470964 580617 471076
rect 580503 470963 580617 470964
rect 581531 410938 581617 485910
rect 582282 473200 582442 503771
rect 583162 496279 583426 504651
rect 583162 496017 583163 496279
rect 583425 496017 583426 496279
rect 583162 496016 583426 496017
rect 583193 488716 583459 488717
rect 583193 488452 583194 488716
rect 583458 488452 583459 488716
rect 583193 488451 583459 488452
rect 582282 473040 582936 473200
rect 582281 472116 582547 472117
rect 582281 471852 582282 472116
rect 582546 471852 582547 472116
rect 582281 471851 582547 471852
rect 581531 410854 581532 410938
rect 581616 410854 581617 410938
rect 581531 410853 581617 410854
rect 582282 407523 582546 471851
rect 582282 407261 582283 407523
rect 582545 407261 582546 407523
rect 582282 407260 582546 407261
rect 505920 390521 506252 390522
rect 480469 390191 505921 390521
rect 506251 390191 506252 390521
rect 505920 390190 506252 390191
rect 451235 389988 451373 389989
rect 77940 389987 451236 389988
rect 77940 389853 77941 389987
rect 78075 389853 451236 389987
rect 77940 389852 451236 389853
rect 451372 389852 451373 389988
rect 451235 389851 451373 389852
rect 450423 389350 450837 389351
rect 78788 389349 450424 389350
rect 78788 388939 78789 389349
rect 79199 388939 450424 389349
rect 78788 388938 450424 388939
rect 450836 388938 450837 389350
rect 450423 388937 450837 388938
rect 449324 388351 449760 388352
rect 79989 388350 449325 388351
rect 79989 388105 79990 388350
rect 80235 388105 449325 388350
rect 79989 388104 449325 388105
rect 302702 387917 449325 388104
rect 449759 387917 449760 388351
rect 449324 387916 449760 387917
rect 442633 387140 443288 387141
rect 72466 386487 442634 387140
rect 443287 386487 443288 387140
rect 72466 386470 72602 386487
rect 442633 386486 443288 386487
rect 439832 385423 439964 385424
rect 71926 385293 439833 385423
rect 439963 385293 439964 385423
rect 439832 385292 439964 385293
rect 441443 384588 442146 384589
rect 71296 383887 441444 384588
rect 442145 383887 442146 384588
rect 441443 383886 442146 383887
rect 439336 383259 439556 383260
rect 70910 383041 439337 383259
rect 439555 383041 439556 383259
rect 16167 376754 16168 376866
rect 16280 376865 69526 376866
rect 16280 376755 69415 376865
rect 69525 376755 69526 376865
rect 16280 376754 69526 376755
rect 16167 376753 16281 376754
rect 70926 349044 71038 383041
rect 439336 383040 439556 383041
rect 438562 382473 438743 382474
rect 71926 382294 438563 382473
rect 438742 382294 438743 382473
rect 71928 352177 72040 382294
rect 438562 382293 438743 382294
rect 90114 381546 158066 381547
rect 90114 381483 158076 381546
rect 90114 381046 150869 381483
rect 150778 380553 150869 381046
rect 157943 380553 158076 381483
rect 150778 380465 158076 380553
rect 128817 380144 132851 380208
rect 128817 380019 128918 380144
rect 90114 379827 128918 380019
rect 132762 380019 132851 380144
rect 132762 379827 132854 380019
rect 90114 379709 132854 379827
rect 136847 379269 140818 379383
rect 136847 379263 136999 379269
rect 90114 378955 136999 379263
rect 136847 378850 136999 378955
rect 140729 379263 140818 379269
rect 140729 378955 140845 379263
rect 140729 378850 140818 378955
rect 136847 378723 140818 378850
rect 128879 377026 132795 377076
rect 128879 376909 128962 377026
rect 72877 376866 72991 376867
rect 90040 376866 128962 376909
rect 72877 376754 72878 376866
rect 72990 376754 128962 376866
rect 72877 376753 72991 376754
rect 90040 376706 128962 376754
rect 128879 376582 128962 376706
rect 132722 376582 132795 377026
rect 128879 376525 132795 376582
rect 417050 371142 440192 380324
rect 545329 376077 548300 376078
rect 452460 376076 545330 376077
rect 452460 373109 452461 376076
rect 455428 373109 545330 376076
rect 452460 373108 545330 373109
rect 548299 373108 548300 376077
rect 545329 373107 548300 373108
rect 90040 369602 158189 369749
rect 90040 366820 150962 369602
rect 157821 366820 158189 369602
rect 90040 366667 158189 366820
rect 90040 364692 132687 364758
rect 90040 363838 128893 364692
rect 132628 363838 132687 364692
rect 90040 363790 132687 363838
rect 90040 362468 140772 362536
rect 90040 361328 136912 362468
rect 140668 361328 140772 362468
rect 90040 361280 140772 361328
rect 71905 352176 72040 352177
rect 71905 352064 71906 352176
rect 72018 352064 72040 352176
rect 71905 352063 72040 352064
rect 71928 352026 72040 352063
rect 82503 356126 130777 356127
rect 82503 355822 130472 356126
rect 130776 355822 130777 356126
rect 82503 355821 130777 355822
rect 13964 348932 71038 349044
rect 13964 334827 14076 348932
rect 15948 345566 16256 345567
rect 82503 345566 82809 355821
rect 15948 345260 15949 345566
rect 16255 345260 82809 345566
rect 83876 354993 139120 354994
rect 83876 354675 138801 354993
rect 139119 354675 139120 354993
rect 83876 354674 139120 354675
rect 15948 345259 16256 345260
rect 15963 344650 16285 344651
rect 83876 344650 84196 354674
rect 15963 344330 15964 344650
rect 16284 344330 84196 344650
rect 90040 347766 169654 352368
rect 90040 345626 116072 347766
rect 118072 345626 169654 347766
rect 15963 344329 16285 344330
rect 15408 343026 83982 343422
rect 90040 343186 169654 345626
rect 15408 339747 15804 343026
rect 16244 342154 82682 342550
rect 15407 339746 15805 339747
rect 15407 339350 15408 339746
rect 15804 339350 15805 339746
rect 15407 339349 15805 339350
rect 16244 338719 16640 342154
rect 25542 341758 81641 341798
rect 25541 341420 81641 341758
rect 25541 340168 26741 341420
rect 27826 340970 77293 341146
rect 27826 340870 28370 340970
rect 28470 340870 77293 340970
rect 27826 340768 77293 340870
rect 27826 340142 29026 340768
rect 16243 338718 16641 338719
rect 16243 338322 16244 338718
rect 16640 338322 16641 338718
rect 16243 338321 16641 338322
rect 76915 337469 77293 340768
rect 81263 338791 81641 341420
rect 82286 339978 82682 342154
rect 83586 341116 83982 343026
rect 83586 340720 154082 341116
rect 82286 339582 109512 339978
rect 159425 338791 159803 343186
rect 81263 338413 159803 338791
rect 76915 337091 109627 337469
rect 44238 334978 44746 334979
rect 13963 334826 14077 334827
rect 13963 334714 13964 334826
rect 14076 334714 14077 334826
rect 13963 334713 14077 334714
rect 44238 334700 44239 334978
rect 42138 334588 44239 334700
rect 14123 333644 14237 333645
rect 14123 333532 14124 333644
rect 14236 333532 14237 333644
rect 14123 333531 14237 333532
rect 14124 325142 14236 333531
rect 42138 325142 42250 334588
rect 44238 334472 44239 334588
rect 44745 334977 131161 334978
rect 44745 334473 130656 334977
rect 131160 334473 131161 334977
rect 44745 334472 131161 334473
rect 44238 334471 44746 334472
rect 44252 334060 44736 334061
rect 44252 333578 44253 334060
rect 44735 334059 139199 334060
rect 44735 333579 138718 334059
rect 139198 333579 139199 334059
rect 44735 333578 139199 333579
rect 44252 333577 44736 333578
rect 14124 325030 42250 325142
rect 86992 314538 114161 314656
rect 86992 311856 106704 314538
rect 113848 311856 114161 314538
rect 86992 311714 114161 311856
rect 86992 310649 132820 310688
rect 86992 310102 128934 310649
rect 132738 310102 132820 310649
rect 86992 310034 132820 310102
rect 86992 309624 140859 309688
rect 86992 309106 136918 309624
rect 140746 309106 140859 309624
rect 86992 309034 140859 309106
rect 15155 307642 15421 307643
rect 15155 307378 15156 307642
rect 15420 307641 17028 307642
rect 15420 307379 16765 307641
rect 17027 307379 17028 307641
rect 15420 307378 17028 307379
rect 15155 307377 15421 307378
rect 13888 302366 14196 302367
rect 13888 302060 13889 302366
rect 14195 302365 130929 302366
rect 14195 302061 130624 302365
rect 130928 302061 130929 302365
rect 14195 302060 130929 302061
rect 13888 302059 14196 302060
rect 14129 301450 14451 301451
rect 14129 301130 14130 301450
rect 14450 301449 138802 301450
rect 14450 301131 138483 301449
rect 138801 301131 138802 301449
rect 14450 301130 138802 301131
rect 14129 301129 14451 301130
rect 13166 297828 153988 298224
rect 13166 296547 13562 297828
rect 13890 297144 109642 297540
rect 13165 296546 13563 296547
rect 13165 296150 13166 296546
rect 13562 296150 13563 296546
rect 13165 296149 13563 296150
rect 13890 295519 14286 297144
rect 32500 295824 32680 295836
rect 32494 295823 32680 295824
rect 32494 295645 32495 295823
rect 32673 295645 32680 295823
rect 13889 295518 14287 295519
rect 13889 295122 13890 295518
rect 14286 295122 14287 295518
rect 32494 295398 32680 295645
rect 13889 295121 14287 295122
rect 31882 294917 32062 294950
rect 31882 294739 31883 294917
rect 32061 294739 32062 294917
rect 14879 281876 15185 281877
rect 14879 281572 14880 281876
rect 15184 281572 15185 281876
rect 14879 259367 15185 281572
rect 15614 281133 15934 281134
rect 15614 280815 15615 281133
rect 15933 280815 15934 281133
rect 14878 259366 15186 259367
rect 14878 259060 14879 259366
rect 15185 259060 15186 259366
rect 14878 259059 15186 259060
rect 15614 258451 15934 280815
rect 31882 274062 32062 294739
rect 32500 274362 32680 295398
rect 100259 286830 169654 290368
rect 66376 285265 67968 285266
rect 100259 285265 122182 286830
rect 66376 283675 66377 285265
rect 67967 284192 122182 285265
rect 124562 284192 169654 286830
rect 292744 286134 292856 352856
rect 435798 349051 438767 371142
rect 577997 349051 580968 349052
rect 435798 346082 577998 349051
rect 580967 346082 580968 349051
rect 577997 346081 580968 346082
rect 582776 321154 582936 473040
rect 583194 451909 583458 488451
rect 583752 479379 583864 479380
rect 583752 479269 583753 479379
rect 583863 479269 583864 479379
rect 583752 457064 583864 479269
rect 583752 457059 583904 457064
rect 583751 457058 583904 457059
rect 583751 456946 583752 457058
rect 583864 456946 583904 457058
rect 583751 456945 583904 456946
rect 583194 451647 583195 451909
rect 583457 451647 583458 451909
rect 583194 451646 583458 451647
rect 583792 450512 583904 456945
rect 583228 450400 583904 450512
rect 583228 412126 583340 450400
rect 583224 412118 583344 412126
rect 583224 412006 583228 412118
rect 583340 412006 583344 412118
rect 583224 412000 583344 412006
rect 582776 320994 583602 321154
rect 582954 319267 583030 319268
rect 582954 319193 582955 319267
rect 583029 319193 583030 319267
rect 571148 318108 571456 318109
rect 453989 318107 571149 318108
rect 453989 317803 453990 318107
rect 454294 317803 571149 318107
rect 453989 317802 571149 317803
rect 571455 317802 571456 318108
rect 571148 317801 571456 317802
rect 571167 317192 571489 317193
rect 446016 317191 571168 317192
rect 446016 316873 446017 317191
rect 446335 316873 571168 317191
rect 446016 316872 571168 316873
rect 571488 316872 571489 317192
rect 571167 316871 571489 316872
rect 582510 315785 582774 315786
rect 582510 315523 582511 315785
rect 582773 315523 582774 315785
rect 571053 312288 571451 312289
rect 432290 311892 571054 312288
rect 571450 311892 571451 312288
rect 571053 311891 571451 311892
rect 419158 310980 448168 311264
rect 571067 311260 571465 311261
rect 419158 310660 444618 310980
rect 419158 301684 419710 310660
rect 423364 301684 444618 310660
rect 419158 301612 444618 301684
rect 447812 301612 448168 310980
rect 469526 310864 469702 311260
rect 470098 310864 571068 311260
rect 571464 310864 571465 311260
rect 571067 310863 571465 310864
rect 582510 310717 582774 315523
rect 582509 310716 582775 310717
rect 582509 310452 582510 310716
rect 582774 310452 582775 310716
rect 582509 310451 582775 310452
rect 419158 301220 448168 301612
rect 305828 299098 456050 299472
rect 305828 299090 452458 299098
rect 305828 292726 306356 299090
rect 313006 292726 452458 299090
rect 305828 292718 452458 292726
rect 455712 292718 456050 299098
rect 305828 292374 456050 292718
rect 417050 287604 477158 290324
rect 67967 283675 169654 284192
rect 66376 283674 67968 283675
rect 66222 281877 66530 281878
rect 66222 281571 66223 281877
rect 66529 281571 93773 281877
rect 66222 281570 66530 281571
rect 66289 281134 66611 281135
rect 66289 280814 66290 281134
rect 66610 280814 92932 281134
rect 66289 280813 66611 280814
rect 77157 279530 77223 279531
rect 77157 279466 77158 279530
rect 77222 279466 77223 279530
rect 77157 279465 77223 279466
rect 77160 278347 77220 279465
rect 92612 278552 92932 280814
rect 93467 279559 93773 281571
rect 100259 281186 169654 283675
rect 417050 284006 427136 287604
rect 430734 284006 477158 287604
rect 417050 283628 477158 284006
rect 477611 283628 477921 283629
rect 417050 283320 477612 283628
rect 477920 283320 477921 283628
rect 417050 281142 477158 283320
rect 477611 283319 477921 283320
rect 93467 279558 131107 279559
rect 93467 279254 130802 279558
rect 131106 279254 131107 279558
rect 93467 279253 131107 279254
rect 571466 278908 571774 278909
rect 453709 278907 571467 278908
rect 453709 278603 453710 278907
rect 454014 278603 571467 278907
rect 453709 278602 571467 278603
rect 571773 278602 571774 278908
rect 571466 278601 571774 278602
rect 92612 278551 138688 278552
rect 77157 278346 77223 278347
rect 77157 278282 77158 278346
rect 77222 278282 77223 278346
rect 77157 278281 77223 278282
rect 92612 278233 138369 278551
rect 138687 278233 138688 278551
rect 92612 278232 138688 278233
rect 571457 277992 571779 277993
rect 446020 277991 571458 277992
rect 66316 277951 67908 277952
rect 66316 276361 66317 277951
rect 67907 276361 91413 277951
rect 446020 277673 446021 277991
rect 446339 277673 571458 277991
rect 446020 277672 571458 277673
rect 571778 277672 571779 277992
rect 571457 277671 571779 277672
rect 66316 276360 67908 276361
rect 89823 275639 91413 276361
rect 582686 276127 582762 276128
rect 582686 276053 582687 276127
rect 582761 276053 582762 276127
rect 32499 274361 32681 274362
rect 32499 274181 32500 274361
rect 32680 274181 32681 274361
rect 32499 274180 32681 274181
rect 31881 274061 32063 274062
rect 31881 273881 31882 274061
rect 32062 273881 32063 274061
rect 89823 274049 109419 275639
rect 31881 273880 32063 273881
rect 571325 273088 571723 273089
rect 430402 272692 571326 273088
rect 571722 272692 571723 273088
rect 571325 272691 571723 272692
rect 571281 272060 571679 272061
rect 469960 271664 571282 272060
rect 571678 271664 571679 272060
rect 571281 271663 571679 271664
rect 563801 261450 563879 261451
rect 582686 261450 582762 276053
rect 563801 261374 563802 261450
rect 563878 261374 582762 261450
rect 563801 261373 563879 261374
rect 15613 258450 15935 258451
rect 15613 258130 15614 258450
rect 15934 258130 15935 258450
rect 15613 258129 15935 258130
rect 563737 256972 563815 256973
rect 582954 256972 583030 319193
rect 583442 276128 583602 320994
rect 583442 276052 583490 276128
rect 583566 276052 583602 276128
rect 583442 276014 583602 276052
rect 563737 256896 563738 256972
rect 563814 256896 583030 256972
rect 583252 274857 583328 274858
rect 583252 274783 583253 274857
rect 583327 274783 583328 274857
rect 563737 256895 563815 256896
rect 466249 255107 473735 255449
rect 563751 255436 563829 255437
rect 583252 255436 583328 274783
rect 563751 255360 563752 255436
rect 563828 255360 583328 255436
rect 563751 255359 563829 255360
rect 15581 253546 15979 253547
rect 15581 253150 15582 253546
rect 15978 253150 15979 253546
rect 15581 253149 15979 253150
rect 14735 252518 15133 252519
rect 14735 252122 14736 252518
rect 15132 252122 15133 252518
rect 14735 252121 15133 252122
rect 11475 247400 11589 247401
rect 11475 247288 11476 247400
rect 11588 247399 13684 247400
rect 11588 247289 13573 247399
rect 13683 247289 13684 247399
rect 11588 247288 13684 247289
rect 11475 247287 11589 247288
rect 14736 222388 15132 252121
rect 15582 223646 15978 253149
rect 466249 247031 466498 255107
rect 473424 252974 473735 255107
rect 477768 252974 478309 252975
rect 473424 252435 477769 252974
rect 478308 252435 478309 252974
rect 473424 247031 473735 252435
rect 477768 252434 478309 252435
rect 476828 247795 525112 247796
rect 476828 247477 476829 247795
rect 477147 247772 525112 247795
rect 477147 247500 524816 247772
rect 525088 247500 525112 247772
rect 477147 247477 525112 247500
rect 476828 247476 525112 247477
rect 462585 245526 462907 245527
rect 453946 245525 462586 245526
rect 453946 245207 453947 245525
rect 454265 245207 462586 245525
rect 453946 245206 462586 245207
rect 462906 245206 462907 245526
rect 462585 245205 462907 245206
rect 462666 244544 463043 244545
rect 445725 244543 462667 244544
rect 445725 244170 445726 244543
rect 446099 244170 462667 244543
rect 445725 244169 462667 244170
rect 463042 244169 463043 244544
rect 462666 244168 463043 244169
rect 103609 234956 130823 234957
rect 103609 234296 130162 234956
rect 130822 234296 130823 234956
rect 103609 234295 130823 234296
rect 69746 224204 70410 224205
rect 103609 224204 104271 234295
rect 15582 223250 23420 223646
rect 69746 223542 69747 224204
rect 70409 223542 104271 224204
rect 105045 233696 139319 233697
rect 105045 233036 138658 233696
rect 139318 233036 139319 233696
rect 105045 233035 139319 233036
rect 69746 223541 70410 223542
rect 69872 223392 70536 223393
rect 105045 223392 105707 233035
rect 69872 222730 69873 223392
rect 70535 222730 105707 223392
rect 106501 232157 114025 232502
rect 106501 224846 106878 232157
rect 113676 224846 114025 232157
rect 69872 222729 70536 222730
rect 106501 222388 114025 224846
rect 14736 221992 114025 222388
rect 4152 220396 9590 220510
rect 4152 215890 4310 220396
rect 9440 215890 9590 220396
rect 4152 215436 9590 215890
rect 4152 210800 4232 215436
rect 9414 210800 9590 215436
rect 4152 210358 9590 210800
rect 4152 205852 4284 210358
rect 9414 205852 9590 210358
rect 4152 205690 9590 205852
rect 106501 201306 114025 221992
rect 466249 221314 473735 247031
rect 574774 240690 580212 240866
rect 574774 236252 574934 240690
rect 580058 236252 580212 240690
rect 574774 235522 580212 236252
rect 574774 231084 574962 235522
rect 580086 231084 580212 235522
rect 574774 230660 580212 231084
rect 574774 226222 574962 230660
rect 580086 226222 580212 230660
rect 574774 226046 580212 226222
rect 466249 211313 466529 221314
rect 473424 211313 473735 221314
rect 466249 210816 473735 211313
rect 106501 194909 106922 201306
rect 113632 194909 114025 201306
rect 106501 194569 114025 194909
rect 574748 196850 580186 197028
rect 574748 192412 574896 196850
rect 580020 192412 580186 196850
rect 574748 192076 580186 192412
rect 451946 191899 580186 192076
rect 451946 187251 452333 191899
rect 455990 187251 580186 191899
rect 451946 187076 580186 187251
rect 574748 186806 580186 187076
rect 532834 185541 533055 185542
rect 532234 185409 532471 185410
rect 531656 185349 531893 185350
rect 531656 185114 531657 185349
rect 531892 185114 531893 185349
rect 444183 180774 448179 180858
rect 444183 179958 444303 180774
rect 448071 180530 448179 180774
rect 448071 180488 475808 180530
rect 448071 180195 479457 180488
rect 448071 180130 475808 180195
rect 448071 179958 448179 180130
rect 444183 179854 448179 179958
rect 3532 178310 8768 178430
rect 3532 173829 3756 178310
rect 8602 173829 8768 178310
rect 452176 177478 456170 177590
rect 452176 176624 452276 177478
rect 456058 177281 456170 177478
rect 456058 177275 475808 177281
rect 456058 176896 478724 177275
rect 456058 176881 475808 176896
rect 456058 176624 456170 176881
rect 452176 176524 456170 176624
rect 3532 173694 8768 173829
rect 466206 175148 473676 175258
rect 3532 173511 133180 173694
rect 3532 168834 129023 173511
rect 132621 168834 133180 173511
rect 466206 173412 466300 175148
rect 473518 174627 473676 175148
rect 473518 173953 477645 174627
rect 473518 173412 473676 173953
rect 466206 173320 473676 173412
rect 3532 168694 133180 168834
rect 3532 168320 8768 168694
rect 3532 163839 3676 168320
rect 8522 163839 8768 168320
rect 3532 163716 8768 163839
rect 417050 167041 475808 170324
rect 417050 163637 431353 167041
rect 434495 163637 475808 167041
rect 417050 161142 475808 163637
rect 89652 146268 169654 150368
rect 474772 148778 475392 161142
rect 476971 149971 477645 173953
rect 478345 150748 478724 176896
rect 479164 151435 479457 180195
rect 510863 151435 511158 151436
rect 479164 151142 510864 151435
rect 511157 151142 511158 151435
rect 510863 151141 511158 151142
rect 511040 150748 511421 150749
rect 478345 150369 511041 150748
rect 511420 150369 511421 150748
rect 511040 150368 511421 150369
rect 510808 149971 511484 149972
rect 476971 149297 510809 149971
rect 511483 149297 511484 149971
rect 510808 149296 511484 149297
rect 511009 148778 511631 148779
rect 474772 148158 511010 148778
rect 511630 148158 511631 148778
rect 511009 148157 511631 148158
rect 89652 143960 146008 146268
rect 148318 143960 169654 146268
rect 89652 141186 169654 143960
rect 22349 136828 130993 136829
rect 22349 136524 130688 136828
rect 130992 136524 130993 136828
rect 22349 136523 130993 136524
rect 22349 131945 22655 136523
rect 23322 136033 139132 136034
rect 23322 135715 138813 136033
rect 139131 135715 139132 136033
rect 23322 135714 139132 135715
rect 22348 131944 22656 131945
rect 22348 131638 22349 131944
rect 22655 131638 22656 131944
rect 22348 131637 22656 131638
rect 23322 131029 23642 135714
rect 78003 133617 79116 133618
rect 144566 133617 145677 141186
rect 78003 132506 78004 133617
rect 79115 132506 145677 133617
rect 78003 132505 79116 132506
rect 78264 131546 78644 131547
rect 78264 131168 78265 131546
rect 78643 131545 130883 131546
rect 78643 131169 130506 131545
rect 130882 131169 130883 131545
rect 78643 131168 130883 131169
rect 78264 131167 78644 131168
rect 23321 131028 23643 131029
rect 23321 130708 23322 131028
rect 23642 130708 23643 131028
rect 23321 130707 23643 130708
rect 78252 129165 78632 129166
rect 78252 128787 78253 129165
rect 78631 129164 139111 129165
rect 78631 128788 138734 129164
rect 139110 128788 139111 129164
rect 78631 128787 139111 128788
rect 78252 128786 78632 128787
rect 47793 127856 48906 127857
rect 47793 126745 47794 127856
rect 48905 126745 109474 127856
rect 47793 126744 48906 126745
rect 23175 126124 23573 126125
rect 23175 125728 23176 126124
rect 23572 125728 153976 126124
rect 23175 125727 23573 125728
rect 23193 125096 23591 125097
rect 23193 124700 23194 125096
rect 23590 124700 110076 125096
rect 23193 124699 23591 124700
rect 77897 119778 78011 119779
rect 77897 119666 77898 119778
rect 78010 119777 130962 119778
rect 78010 119667 130809 119777
rect 130919 119667 130962 119777
rect 78010 119666 130962 119667
rect 77897 119665 78011 119666
rect 128818 119218 280542 119470
rect 128818 112664 129090 119218
rect 132624 119060 280542 119218
rect 132624 112664 273522 119060
rect 128818 112606 273522 112664
rect 280172 112606 280542 119060
rect 128818 112302 280542 112606
rect 444175 92247 448174 92351
rect 444175 91356 444290 92247
rect 448055 92019 448174 92247
rect 448055 91619 480762 92019
rect 448055 91356 448174 91619
rect 444175 91248 448174 91356
rect 452177 89388 456180 89459
rect 452177 89142 452241 89388
rect 29440 88744 29748 88745
rect 29440 88438 29441 88744
rect 29747 88743 130975 88744
rect 29747 88439 130670 88743
rect 130974 88439 130975 88743
rect 452171 88742 452241 89142
rect 29747 88438 130975 88439
rect 452177 88492 452241 88742
rect 456105 89142 456180 89388
rect 456105 88742 480762 89142
rect 456105 88492 456180 88742
rect 29440 88437 29748 88438
rect 452177 88434 456180 88492
rect 29645 87828 29967 87829
rect 29645 87508 29646 87828
rect 29966 87827 139272 87828
rect 29966 87509 138953 87827
rect 139271 87509 139272 87827
rect 29966 87508 139272 87509
rect 29645 87507 29967 87508
rect 29595 82924 29993 82925
rect 29595 82528 29596 82924
rect 29992 82528 154456 82924
rect 29595 82527 29993 82528
rect 29603 81896 30001 81897
rect 29603 81500 29604 81896
rect 30000 81500 109984 81896
rect 29603 81499 30001 81500
rect 120565 81344 120963 81345
rect 120565 80948 120566 81344
rect 120962 80948 154356 81344
rect 120565 80947 120963 80948
rect 446266 74825 503305 74826
rect 446266 74534 446267 74825
rect 446558 74534 503305 74825
rect 446266 74533 503305 74534
rect 453465 73948 502642 73949
rect 453465 73571 453466 73948
rect 453843 73571 502642 73948
rect 453465 73570 502642 73571
rect 39720 71358 146167 72920
rect 468962 71497 469417 72171
rect 470091 71497 501577 72171
rect 144605 67029 146167 71358
rect 150028 67029 169654 70368
rect 144605 66158 169654 67029
rect 144605 65467 159964 66158
rect 150028 63802 159964 65467
rect 162104 63802 169654 66158
rect 150028 61186 169654 63802
rect 417050 67289 480762 70324
rect 417050 63691 436136 67289
rect 439734 64614 480762 67289
rect 439734 63994 500184 64614
rect 439734 63691 480762 63994
rect 417050 61142 480762 63691
rect 42785 59527 139161 59528
rect 42785 58139 42786 59527
rect 44174 58139 137772 59527
rect 139160 58139 139161 59527
rect 42785 58138 139161 58139
rect 466219 59292 473683 59375
rect 466219 58179 466321 59292
rect 473542 58976 473683 59292
rect 473542 58576 480762 58976
rect 473542 58179 473683 58576
rect 466219 58099 473683 58179
rect 499564 52876 500184 63994
rect 500903 54009 501577 71497
rect 502263 54732 502642 73570
rect 503012 55249 503305 74533
rect 531656 63772 531893 185114
rect 532234 185174 532235 185409
rect 532470 185174 532471 185409
rect 532234 161950 532471 185174
rect 532834 185322 532835 185541
rect 533054 185322 533055 185541
rect 532233 161949 532472 161950
rect 532233 161712 532234 161949
rect 532471 161712 532472 161949
rect 532233 161711 532472 161712
rect 531655 63771 531894 63772
rect 531655 63534 531656 63771
rect 531893 63534 531894 63771
rect 531655 63533 531894 63534
rect 527285 55249 527580 55250
rect 503012 54956 527286 55249
rect 527579 54956 527580 55249
rect 527285 54955 527580 54956
rect 527332 54732 527713 54733
rect 502263 54353 527333 54732
rect 527712 54353 527713 54732
rect 527332 54352 527713 54353
rect 527694 54009 528370 54010
rect 500903 53335 527695 54009
rect 528369 53335 528370 54009
rect 527694 53334 528370 53335
rect 527851 52876 528473 52877
rect 499564 52256 527852 52876
rect 528472 52256 528473 52876
rect 527851 52255 528473 52256
rect 39800 46645 131774 46646
rect 24124 45544 24432 45545
rect 24124 45238 24125 45544
rect 24431 45238 28889 45544
rect 24124 45237 24432 45238
rect 24085 44628 24407 44629
rect 24085 44308 24086 44628
rect 24406 44308 27940 44628
rect 24085 44307 24407 44308
rect 27620 43224 27940 44308
rect 28583 44077 28889 45238
rect 39800 45059 130143 46645
rect 131729 45059 131774 46645
rect 39800 45058 131774 45059
rect 28583 44076 130967 44077
rect 28583 43772 130662 44076
rect 130966 43772 130967 44076
rect 28583 43771 130967 43772
rect 27620 43223 138916 43224
rect 27620 42905 138597 43223
rect 138915 42905 138916 43223
rect 27620 42904 138916 42905
rect 102396 41327 120962 41328
rect 102396 40933 120567 41327
rect 120961 40933 120962 41327
rect 102396 40932 120962 40933
rect 23431 39724 23829 39725
rect 102396 39724 102792 40932
rect 23431 39328 23432 39724
rect 23828 39328 102792 39724
rect 136362 40865 167859 41116
rect 23431 39327 23829 39328
rect 106528 38790 114018 38902
rect 23401 38696 23799 38697
rect 106528 38696 106610 38790
rect 23401 38300 23402 38696
rect 23798 38300 106610 38696
rect 23401 38299 23799 38300
rect 106528 38256 106610 38300
rect 113894 38696 114018 38790
rect 113894 38300 114056 38696
rect 113894 38256 114018 38300
rect 106528 38162 114018 38256
rect 136362 31547 137083 40865
rect 140503 31610 157632 40865
rect 167451 31610 167859 40865
rect 426799 39173 434047 39338
rect 426799 32240 426979 39173
rect 433851 32240 434047 39173
rect 426799 32090 434047 32240
rect 140503 31547 167859 31610
rect 136362 31139 167859 31547
rect 531656 23016 531893 63533
rect 532234 49008 532471 161711
rect 532834 81407 533055 185322
rect 574748 182368 574908 186806
rect 580032 182368 580186 186806
rect 574748 182208 580186 182368
rect 533413 179627 533636 179628
rect 533413 179406 533414 179627
rect 533635 179406 533636 179627
rect 533413 179405 533636 179406
rect 533414 93713 533635 179405
rect 551028 148777 551648 155236
rect 551028 148159 551029 148777
rect 551647 148159 551648 148777
rect 551028 148158 551648 148159
rect 574794 152256 580634 152400
rect 574794 147818 575156 152256
rect 580280 147818 580634 152256
rect 574794 147254 580634 147818
rect 574794 142816 575132 147254
rect 580256 142816 580634 147254
rect 574794 142194 580634 142816
rect 574794 137756 575102 142194
rect 580226 137756 580634 142194
rect 574794 137630 580634 137756
rect 533414 93712 560748 93713
rect 533414 93493 560528 93712
rect 560747 93493 560748 93712
rect 533414 93492 560748 93493
rect 532833 81406 533056 81407
rect 532833 81185 532834 81406
rect 533055 81185 533056 81406
rect 532833 81184 533056 81185
rect 532234 48896 532272 49008
rect 532384 48896 532471 49008
rect 532234 48794 532471 48896
rect 532834 25352 533055 81184
rect 552580 52875 553200 57058
rect 552580 52257 552581 52875
rect 553199 52257 553200 52875
rect 552580 52256 553200 52257
rect 3527 18189 460533 18190
rect 3527 18157 124736 18189
rect 3527 17264 3562 18157
rect 4344 17264 124736 18157
rect 3527 17233 124736 17264
rect 125692 17233 459576 18189
rect 460532 17233 460533 18189
rect 531698 17823 531810 23016
rect 532878 22551 532990 25352
rect 532877 22550 532991 22551
rect 532877 22438 532878 22550
rect 532990 22438 532991 22550
rect 532877 22437 532991 22438
rect 531697 17822 531811 17823
rect 531697 17710 531698 17822
rect 531810 17710 531811 17822
rect 531697 17709 531811 17710
rect 3527 17232 460533 17233
<< via4 >>
rect 516456 693856 520966 698932
rect 107279 598134 108964 599819
rect 107507 586760 109192 588445
rect 469329 595339 471323 597333
rect 430382 586892 430778 587288
rect 469412 585864 469808 586260
rect 107787 579654 109472 581339
rect 108171 568273 109856 569958
rect 4066 555362 9170 560048
rect 466599 553646 473439 560021
rect 575622 546532 580746 550970
rect 466547 523885 473413 530621
rect 154256 518376 154652 518772
rect 109858 517542 110254 517938
rect 469384 505064 469780 505460
rect 430442 503372 430838 503768
rect 109971 497730 110368 498127
rect 429948 491342 430344 491738
rect 469798 490244 470194 490640
rect 469678 488997 470107 489426
rect 430200 480314 430596 480710
rect 154442 479222 154838 479618
rect 470294 479056 470690 479452
rect 106611 470309 113894 475380
rect 273502 472070 280420 478254
rect 150899 461395 157916 462824
rect 106619 454319 113903 455661
rect 106630 440408 113902 441575
rect 150941 439040 157881 440395
rect 153732 434810 154128 435206
rect 109890 434164 110286 434560
rect 154300 402698 154696 403094
rect 109920 391468 110316 391864
rect 163821 391614 167356 400684
rect 150869 380553 157943 381483
rect 150962 366820 157821 369602
rect 154082 340720 154478 341116
rect 109512 339582 109908 339978
rect 109627 337091 110005 337469
rect 106704 311856 113848 314538
rect 153988 297828 154384 298224
rect 109642 297144 110038 297540
rect 431894 311892 432290 312288
rect 419710 301684 423364 310660
rect 469702 310864 470098 311260
rect 306356 292726 313006 299090
rect 109419 274049 111009 275639
rect 430006 272692 430402 273088
rect 469564 271664 469960 272060
rect 466498 247031 473424 255107
rect 524816 247500 525088 247772
rect 23420 223250 23816 223646
rect 106878 224846 113676 232157
rect 4232 210800 9414 215436
rect 574962 231084 580086 235522
rect 466529 211313 473424 221314
rect 106922 194909 113632 201306
rect 466300 173412 473518 175148
rect 109474 126745 110585 127856
rect 153976 125728 154372 126124
rect 110076 124700 110472 125096
rect 273522 112606 280172 119060
rect 154456 82528 154852 82924
rect 109984 81500 110380 81896
rect 154356 80948 154752 81344
rect 469417 71497 470091 72171
rect 466321 58179 473542 59292
rect 106610 38256 113894 38790
rect 157632 31610 167451 40865
rect 426979 32240 433851 39173
rect 575132 142816 580256 147254
<< metal5 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 516238 698932 521238 699090
rect 516238 696670 516456 698932
rect 515321 693856 516456 696670
rect 520966 696670 521238 698932
rect 520966 693856 522787 696670
rect 515321 672866 522787 693856
rect 106520 665257 280703 672722
rect 106520 599819 114019 665257
rect 106520 598134 107279 599819
rect 108964 598134 114019 599819
rect 106520 588445 114019 598134
rect 106520 586760 107507 588445
rect 109192 586760 114019 588445
rect 106520 581339 114019 586760
rect 106520 579654 107787 581339
rect 109472 579654 114019 581339
rect 106520 569958 114019 579654
rect 106520 568273 108171 569958
rect 109856 568273 114019 569958
rect 106520 561595 114019 568273
rect 6412 560186 114019 561595
rect 3942 560048 114019 560186
rect 3942 555362 4066 560048
rect 9170 555362 114019 560048
rect 3942 555186 114019 555362
rect 6412 554130 114019 555186
rect 106520 517938 114019 554130
rect 106520 517542 109858 517938
rect 110254 517542 114019 517938
rect 106520 498127 114019 517542
rect 106520 497730 109971 498127
rect 110368 497730 114019 498127
rect 106520 475380 114019 497730
rect 106520 470309 106611 475380
rect 113894 470309 114019 475380
rect 106520 455661 114019 470309
rect 106520 454319 106619 455661
rect 113903 454319 114019 455661
rect 106520 441575 114019 454319
rect 106520 440408 106630 441575
rect 113902 440408 114019 441575
rect 106520 434560 114019 440408
rect 106520 434164 109890 434560
rect 110286 434164 114019 434560
rect 106520 391864 114019 434164
rect 106520 391468 109920 391864
rect 110316 391468 114019 391864
rect 106520 339978 114019 391468
rect 106520 339582 109512 339978
rect 109908 339582 114019 339978
rect 106520 337469 114019 339582
rect 106520 337091 109627 337469
rect 110005 337091 114019 337469
rect 106520 314538 114019 337091
rect 106520 311856 106704 314538
rect 113848 311856 114019 314538
rect 106520 297540 114019 311856
rect 106520 297144 109642 297540
rect 110038 297144 114019 297540
rect 106520 275639 114019 297144
rect 106520 274049 109419 275639
rect 111009 274049 114019 275639
rect 106520 232157 114019 274049
rect 106520 224846 106878 232157
rect 113676 224846 114019 232157
rect 106520 224434 114019 224846
rect 150783 572691 172377 579941
rect 150783 518772 158033 572691
rect 150783 518376 154256 518772
rect 154652 518376 158033 518772
rect 150783 489095 158033 518376
rect 273238 490588 280703 665257
rect 305969 665400 522787 672866
rect 150783 481845 169318 489095
rect 273238 483123 292180 490588
rect 273238 483118 280703 483123
rect 150783 479618 158033 481845
rect 150783 479222 154442 479618
rect 154838 479222 158033 479618
rect 150783 462824 158033 479222
rect 150783 461395 150899 462824
rect 157916 461395 158033 462824
rect 150783 440395 158033 461395
rect 150783 439040 150941 440395
rect 157881 439040 158033 440395
rect 150783 435206 158033 439040
rect 150783 434810 153732 435206
rect 154128 434810 158033 435206
rect 150783 403094 158033 434810
rect 150783 402698 154300 403094
rect 154696 402698 158033 403094
rect 150783 381483 158033 402698
rect 273238 478254 280703 479132
rect 273238 472070 273502 478254
rect 280420 472070 280703 478254
rect 163332 400684 168774 401219
rect 163332 391614 163821 400684
rect 167356 391614 168774 400684
rect 163332 391172 168774 391614
rect 273238 388006 280703 472070
rect 284715 382048 292180 483123
rect 305969 400556 313435 665400
rect 466215 597333 473681 665400
rect 466215 595339 469329 597333
rect 471323 595339 473681 597333
rect 426804 587288 434054 590775
rect 426804 586892 430382 587288
rect 430778 586892 434054 587288
rect 426804 579339 434054 586892
rect 418431 572089 434054 579339
rect 426804 546276 434054 572089
rect 466215 586260 473681 595339
rect 466215 585864 469412 586260
rect 469808 585864 473681 586260
rect 466215 560021 473681 585864
rect 466215 553646 466599 560021
rect 473439 553646 473681 560021
rect 466215 553211 473681 553646
rect 553960 551280 577018 551988
rect 553960 550970 580932 551280
rect 553960 546532 575622 550970
rect 580746 546532 580932 550970
rect 553960 546280 580932 546532
rect 553960 546276 577018 546280
rect 426804 544738 577018 546276
rect 426804 539026 561210 544738
rect 426804 503768 434054 539026
rect 426804 503372 430442 503768
rect 430838 503372 434054 503768
rect 426804 491738 434054 503372
rect 426804 491342 429948 491738
rect 430344 491342 434054 491738
rect 426804 489339 434054 491342
rect 418431 482089 434054 489339
rect 426804 480710 434054 482089
rect 426804 480314 430200 480710
rect 430596 480314 434054 480710
rect 426804 430706 434054 480314
rect 426216 427736 434054 430706
rect 150783 380553 150869 381483
rect 157943 380553 158033 381483
rect 150783 369602 158033 380553
rect 150783 366820 150962 369602
rect 157821 366820 158033 369602
rect 150783 341116 158033 366820
rect 150783 340720 154082 341116
rect 154478 340720 158033 341116
rect 150783 309095 158033 340720
rect 273238 374583 292180 382048
rect 295875 393090 313435 400556
rect 426804 399339 434054 427736
rect 466215 530621 473681 530943
rect 466215 523885 466547 530621
rect 473413 523885 473681 530621
rect 466215 505460 473681 523885
rect 466215 505064 469384 505460
rect 469780 505064 473681 505460
rect 466215 490640 473681 505064
rect 466215 490244 469798 490640
rect 470194 490244 473681 490640
rect 466215 489426 473681 490244
rect 466215 488997 469678 489426
rect 470107 488997 473681 489426
rect 466215 479452 473681 488997
rect 466215 479056 470294 479452
rect 470690 479056 473681 479452
rect 466215 412769 473681 479056
rect 466206 409865 473703 412769
rect 150783 301845 169318 309095
rect 150783 298224 158033 301845
rect 150783 297828 153988 298224
rect 154384 297828 158033 298224
rect 23396 223646 23840 223670
rect 23396 223250 23420 223646
rect 23816 223250 23840 223646
rect 23396 223226 23840 223250
rect 23420 216733 23816 223226
rect 150783 219095 158033 297828
rect 150783 216733 169318 219095
rect 8595 215634 169318 216733
rect 4098 215436 169318 215634
rect 4098 210800 4232 215436
rect 9414 211845 169318 215436
rect 9414 210800 158033 211845
rect 4098 210634 158033 210800
rect 8595 209483 158033 210634
rect 106520 201306 114019 201663
rect 106520 194909 106922 201306
rect 113632 194909 114019 201306
rect 106520 127856 114019 194909
rect 106520 126745 109474 127856
rect 110585 126745 114019 127856
rect 106520 125096 114019 126745
rect 106520 124700 110076 125096
rect 110472 124700 114019 125096
rect 106520 81896 114019 124700
rect 106520 81500 109984 81896
rect 110380 81500 114019 81896
rect 106520 38790 114019 81500
rect 150783 129095 158033 209483
rect 150783 126124 169318 129095
rect 150783 125728 153976 126124
rect 154372 125728 169318 126124
rect 150783 121845 169318 125728
rect 273238 123226 280703 374583
rect 295875 289002 303341 393090
rect 418431 392089 434054 399339
rect 305969 299090 313435 378716
rect 426804 312288 434054 392089
rect 426804 311892 431894 312288
rect 432290 311892 434054 312288
rect 418572 310660 423932 311208
rect 418572 301684 419710 310660
rect 423364 301684 423932 310660
rect 426804 309339 434054 311892
rect 426752 302089 434054 309339
rect 418572 301208 423932 301684
rect 305969 292726 306356 299090
rect 313006 292726 313435 299090
rect 305969 291859 313435 292726
rect 295875 289000 313304 289002
rect 295875 281529 313435 289000
rect 150783 82924 158033 121845
rect 150783 82528 154456 82924
rect 154852 82528 158033 82924
rect 150783 81344 158033 82528
rect 150783 80948 154356 81344
rect 154752 80948 158033 81344
rect 150783 77477 158033 80948
rect 273238 119060 280703 119494
rect 273238 112606 273522 119060
rect 280172 112606 280703 119060
rect 106520 38256 106610 38790
rect 113894 38256 114019 38790
rect 106520 38157 114019 38256
rect 157255 40865 168455 41208
rect 157255 31610 157632 40865
rect 167451 31610 168455 40865
rect 157255 31208 168455 31610
rect 273238 31207 280703 112606
rect 305969 26129 313435 281529
rect 426804 273088 434054 302089
rect 426804 272692 430006 273088
rect 430402 272692 434054 273088
rect 426804 237151 434054 272692
rect 466215 368506 473681 409865
rect 466215 366922 473688 368506
rect 466215 311260 473681 366922
rect 466215 310864 469702 311260
rect 470098 310864 473681 311260
rect 466215 272060 473681 310864
rect 466215 271664 469564 272060
rect 469960 271664 473681 272060
rect 466215 255107 473681 271664
rect 466215 247031 466498 255107
rect 473424 247031 473681 255107
rect 524792 247772 526584 247796
rect 524792 247500 524816 247772
rect 525088 247500 526584 247772
rect 524792 247476 526584 247500
rect 466215 246663 473681 247031
rect 426804 235850 577018 237151
rect 426804 235522 580166 235850
rect 426804 231084 574962 235522
rect 580086 231084 580166 235522
rect 426804 230850 580166 231084
rect 426804 229901 577018 230850
rect 426804 219339 434054 229901
rect 418431 212089 434054 219339
rect 426804 129339 434054 212089
rect 418431 122089 434054 129339
rect 426804 39339 434054 122089
rect 418431 39173 434054 39339
rect 418431 32240 426979 39173
rect 433851 32240 434054 39173
rect 418431 32089 434054 32240
rect 466215 221314 473681 221672
rect 466215 211313 466529 221314
rect 473424 211313 473681 221314
rect 466215 175148 473681 211313
rect 466215 173412 466300 175148
rect 473518 173412 473681 175148
rect 466215 103777 473681 173412
rect 573526 149883 580992 153349
rect 573534 147254 580992 149883
rect 573534 142816 575132 147254
rect 580256 142816 580992 147254
rect 573534 139533 580992 142816
rect 573526 103777 580992 139533
rect 466215 96311 580992 103777
rect 466215 72171 473681 96311
rect 466215 71497 469417 72171
rect 470091 71497 473681 72171
rect 466215 59292 473681 71497
rect 466215 58179 466321 59292
rect 473542 58179 473681 59292
rect 466215 26129 473681 58179
rect 305969 18663 473687 26129
<< fillblock >>
rect 287497 306699 302657 310031
rect 290225 302778 296473 306103
<< comment >>
rect 0 704800 585600 705600
rect 0 800 800 704800
rect 584800 800 585600 704800
rect 0 0 585600 800
use ct2_switch_array  ct2_switch_array_0
timestamp 1726321856
transform 1 0 -186 0 1 84470
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_1
timestamp 1726321856
transform 1 0 378 0 1 -215552
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_2
timestamp 1726321856
transform 1 0 -186 0 1 41270
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_3
timestamp 1726321856
transform 1 0 -186 0 1 127870
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_4
timestamp 1726321856
transform 1 0 -186 0 1 171070
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_5
timestamp 1726321856
transform 1 0 -186 0 1 214270
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_6
timestamp 1726321856
transform 1 0 -186 0 1 257470
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_7
timestamp 1726321856
transform 1 0 -186 0 1 -1730
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_8
timestamp 1726321856
transform 1 0 378 0 1 -129152
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_9
timestamp 1726321856
transform 1 0 378 0 1 -172352
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_10
timestamp 1726321856
transform -1 0 584704 0 1 332012
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_11
timestamp 1726321856
transform -1 0 584704 0 1 17812
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_12
timestamp 1726321856
transform -1 0 584704 0 1 57012
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_13
timestamp 1726321856
transform -1 0 584704 0 1 218412
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_14
timestamp 1726321856
transform -1 0 584704 0 1 251212
box 2132 252898 13728 266392
use ct2_switch_array  ct2_switch_array_15
timestamp 1726321856
transform -1 0 584704 0 1 235012
box 2132 252898 13728 266392
use font_4C  font_4C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766404
transform 1 0 295208 0 1 507055
box 0 0 1080 2520
use font_4F  font_4F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598767855
transform 1 0 296660 0 1 507074
box 0 0 1080 2520
use font_4F  font_4F_1
timestamp 1598767855
transform 1 0 298113 0 1 507092
box 0 0 1080 2520
use font_5A  font_5A_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598772956
transform 1 0 299565 0 1 507111
box 0 0 1080 2520
use font_30  font_30_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786981
transform 1 0 292120 0 1 503139
box 0 0 1080 2520
use font_32  font_32_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787041
transform 1 0 290686 0 1 503118
box 0 0 1080 2520
use font_32  font_32_1
timestamp 1598787041
transform 1 0 293535 0 1 503118
box 0 0 1080 2520
use font_34  font_34_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787136
transform 1 0 295024 0 1 503154
box 0 0 1080 2520
use font_41  font_41_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763107
transform 1 0 293756 0 1 507074
box 0 0 1080 2520
use font_41  font_41_1
timestamp 1598763107
transform 1 0 300982 0 1 507129
box 0 0 1080 2520
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 287836 0 1 507088
box 0 0 1080 2520
use font_48  font_48_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765560
transform 1 0 289326 0 1 507111
box 0 0 1080 2520
use font_49  font_49_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765816
transform 1 0 290833 0 1 507111
box 0 0 1080 2520
use font_50  font_50_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 292285 0 1 507092
box 0 0 1080 2520
use power_stage  power_stage_0 ../dependencies/sky130_ef_ip__analog_switches/mag
array 0 6 90000 0 0 -111006
timestamp 1714671808
transform 0 -1 234941 1 0 120408
box -89200 -44204 -9499 66802
use power_stage  power_stage_1
array 0 6 90000 0 0 111006
timestamp 1714671808
transform 0 1 351850 1 0 120408
box -89200 -44204 -9499 66802
use sky130_aa_ip__programmable_pll  sky130_aa_ip__programmable_pll_0 ../dependencies/sky130_aa_ip__programmable_pll/mag
timestamp 1726362604
transform 1 0 482169 0 1 380775
box -34505 -65703 98798 121313
use sky130_ak_ip__cmos_vref  sky130_ak_ip__cmos_vref_0 ../dependencies/sky130_ak_ip__cmos_vref/mag
timestamp 1721067183
transform -1 0 61111 0 1 433301
box 8587 -19903 21921 206
use sky130_am_ip__ldo_01v8  sky130_am_ip__ldo_01v8_0 ../dependencies/sky130_am_ip__ldo_01v8/mag
timestamp 1721052427
transform 0 -1 40439 1 0 487967
box 4253 -10775 28439 6899
use sky130_ef_ip__ccomp3v_cl  sky130_ef_ip__ccomp3v_cl_0 ../dependencies/sky130_ef_ip__ccomp3v/mag
timestamp 1721179627
transform 1 0 25256 0 1 330161
box -322 -2743 13304 10357
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../dependencies/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1724445404
transform -1 0 114444 0 -1 238850
box 52849 -36868 89580 14592
use sky130_ef_ip__idac3v_8bit  sky130_ef_ip__idac3v_8bit_0 ../dependencies/sky130_ef_ip__biasgen/mag
timestamp 1724460830
transform -1 0 73100 0 -1 601014
box -1186 -1691 49914 35112
use sky130_ef_ip__rc_osc_16M  sky130_ef_ip__rc_osc_16M_0 ../dependencies/sky130_ef_ip__rc_osc_16M/mag
timestamp 1721245376
transform 1 0 30916 0 1 124804
box 0 700 10977 10024
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_1 ../dependencies/sky130_ef_ip__rc_osc_500k/mag
timestamp 1721241604
transform 1 0 546532 0 1 605912
box 0 0 12242 10724
use sky130_ef_ip__rdac3v_8bit  sky130_ef_ip__rdac3v_8bit_0 ../dependencies/sky130_ef_ip__rdac3v_8bit/mag
timestamp 1718228761
transform 0 1 536300 1 0 56638
box -200 -200 25939 21270
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_0 ../dependencies/sky130_ef_ip__rheostat_8bit/mag
timestamp 1716082924
transform 0 1 534748 1 0 154816
box -200 -4 25939 16904
use sky130_ef_ip__samplehold  sky130_ef_ip__samplehold_0 ../dependencies/sky130_ef_ip__samplehold/mag
timestamp 1718244471
transform 1 0 533435 0 1 513311
box 537 303 14883 11558
use sky130_icrg_ip__ulpcomp2  sky130_icrg_ip__ulpcomp2_0 ../dependencies/sky130_icrg_ip__ulpcomp/mag
timestamp 1720377809
transform 1 0 533375 0 -1 481444
box -625 -8056 8504 1566
use sky130_iic_ip__audiodac_drv_lite  sky130_iic_ip__audiodac_drv_lite_0 ../dependencies/sky130_iic_ip__audiodac_v1/mag
timestamp 1724508986
transform -1 0 40116 0 1 44674
box -316 -300 9632 28678
use sky130_sw_ip__bgrref_por  sky130_sw_ip__bgrref_por_0 ../dependencies/sky130_sw_ip__bgrref_por/mag
timestamp 1721440821
transform 1 0 523787 0 1 545780
box 2359 -300396 39662 -277894
<< labels >>
flabel metal4 15162 171077 15162 171077 0 FreeSans 16000 0 0 0 vssd2
flabel metal4 13496 642110 13496 642110 0 FreeSans 16000 0 0 0 vccd2
flabel metal2 s 180988 0 181100 1280 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 184534 0 184646 1280 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 195172 0 195284 1280 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 198718 0 198830 1280 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 202264 0 202376 1280 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205810 0 205922 1280 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 209356 0 209468 1280 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 216448 0 216560 1280 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219994 0 220106 1280 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 223540 0 223652 1280 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 227086 0 227198 1280 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 230632 0 230744 1280 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 234178 0 234290 1280 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 237724 0 237836 1280 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 241270 0 241382 1280 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244816 0 244928 1280 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 248362 0 248474 1280 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251908 0 252020 1280 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 255454 0 255566 1280 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 259000 0 259112 1280 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 262546 0 262658 1280 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 266092 0 266204 1280 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 269638 0 269750 1280 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 273184 0 273296 1280 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 276730 0 276842 1280 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 280276 0 280388 1280 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283822 0 283934 1280 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 287368 0 287480 1280 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290914 0 291026 1280 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 294460 0 294572 1280 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 298006 0 298118 1280 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 301552 0 301664 1280 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 305098 0 305210 1280 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 308644 0 308756 1280 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 312190 0 312302 1280 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 315736 0 315848 1280 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 319282 0 319394 1280 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322828 0 322940 1280 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 326374 0 326486 1280 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329920 0 330032 1280 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 333466 0 333578 1280 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 337012 0 337124 1280 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 340558 0 340670 1280 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 344104 0 344216 1280 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 347650 0 347762 1280 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 351196 0 351308 1280 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 354742 0 354854 1280 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 358288 0 358400 1280 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361834 0 361946 1280 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 365380 0 365492 1280 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368926 0 369038 1280 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 372472 0 372584 1280 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 376018 0 376130 1280 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 379564 0 379676 1280 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 383110 0 383222 1280 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 386656 0 386768 1280 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 390202 0 390314 1280 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 393748 0 393860 1280 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 397294 0 397406 1280 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400840 0 400952 1280 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 404386 0 404498 1280 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407932 0 408044 1280 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 411478 0 411590 1280 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 415024 0 415136 1280 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 418570 0 418682 1280 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 422116 0 422228 1280 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 425662 0 425774 1280 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 429208 0 429320 1280 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 432754 0 432866 1280 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 436300 0 436412 1280 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439846 0 439958 1280 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 443392 0 443504 1280 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 446938 0 447050 1280 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 450484 0 450596 1280 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 454030 0 454142 1280 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 457576 0 457688 1280 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 461122 0 461234 1280 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 464668 0 464780 1280 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 468214 0 468326 1280 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 471760 0 471872 1280 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 475306 0 475418 1280 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478852 0 478964 1280 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 482398 0 482510 1280 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485944 0 486056 1280 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 489490 0 489602 1280 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 493036 0 493148 1280 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 496582 0 496694 1280 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 500128 0 500240 1280 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 503674 0 503786 1280 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 507220 0 507332 1280 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 510766 0 510878 1280 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 514312 0 514424 1280 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 517858 0 517970 1280 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 521404 0 521516 1280 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524950 0 525062 1280 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 528496 0 528608 1280 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 532042 0 532154 1280 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 535588 0 535700 1280 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 539134 0 539246 1280 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541498 0 541610 1280 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 545044 0 545156 1280 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 548590 0 548702 1280 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 552136 0 552248 1280 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 556864 0 556976 1280 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 560410 0 560522 1280 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563956 0 564068 1280 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 567502 0 567614 1280 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal3 s 583100 678784 585600 683784 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 584320 590272 585600 590384 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s 584320 589090 585600 589202 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s 584320 584362 585600 584474 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 584320 500850 585600 500962 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 584320 499668 585600 499780 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 584320 494940 585600 495052 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 584320 451700 585600 451812 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 584320 407278 585600 407390 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 584320 360856 585600 360968 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 584320 314452 585600 314564 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 584320 275940 585600 276052 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 584320 274758 585600 274870 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 584320 270030 585600 270142 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s 584320 95918 585600 96030 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 584320 94736 585600 94848 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 584320 51260 585600 51372 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 584320 50078 585600 50190 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 584320 24802 585600 24914 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 584320 23620 585600 23732 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 584320 20074 585600 20186 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 584320 18892 585600 19004 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 584320 15346 585600 15458 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 584320 14164 585600 14276 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 584320 10618 585600 10730 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s 584320 9436 585600 9548 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s 584320 5890 585600 6002 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 584320 320362 585600 320474 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 584320 319180 585600 319292 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 584320 4708 585600 4820 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 800 163688 2460 168488 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal3 s 800 550242 2460 555042 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 800 205688 2460 210488 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 800 634642 2460 639442 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 567394 703100 572394 705600 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 521394 703140 526194 705600 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 511394 703140 516194 705600 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 466194 703100 471194 705600 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 414194 703100 419194 705600 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 330094 703100 335094 705600 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 218094 703100 223094 705600 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 166394 703100 171394 705600 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 120994 703100 125994 705600 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68994 703100 73994 705600 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16994 703100 21994 705600 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 800 681042 2500 686042 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 800 644642 2460 649442 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 800 560242 2460 565042 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 511148 1280 511260 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s 0 469108 1280 469220 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s 0 425886 1280 425998 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 0 382664 1280 382776 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 0 377936 1280 378048 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s 0 376754 1280 376866 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s 0 339442 1280 339554 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s 0 296220 1280 296332 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s 0 253198 1280 253310 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s 800 215688 2460 220488 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 800 173688 2460 178488 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 125576 1280 125688 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s 0 82354 1280 82466 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s 0 39132 1280 39244 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s 0 34404 1280 34516 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s 0 33222 1280 33334 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s 0 17710 1280 17822 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 0 12982 1280 13094 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s 0 11800 1280 11912 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s 0 8254 1280 8366 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s 0 7072 1280 7184 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s 583140 137630 585600 142430 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 583140 182230 585600 187030 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 583140 226030 585600 230830 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 583140 541362 585600 546162 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 583140 630584 585600 635384 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal2 s 571048 0 571160 1280 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 191626 0 191738 1280 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 188080 0 188192 1280 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 131344 0 131456 1280 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 134890 0 135002 1280 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 138436 0 138548 1280 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 141982 0 142094 1280 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 145528 0 145640 1280 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 149074 0 149186 1280 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 152620 0 152732 1280 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 156166 0 156278 1280 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 159712 0 159824 1280 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 163258 0 163370 1280 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 166804 0 166916 1280 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 170350 0 170462 1280 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173896 0 174008 1280 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 177442 0 177554 1280 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal4 42979 17673 42979 17673 0 FreeSans 16000 0 0 0 bias_reference_voltage
<< end >>
